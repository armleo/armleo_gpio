VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO armleo_gpio
  CLASS BLOCK ;
  FOREIGN armleo_gpio ;
  ORIGIN 0.000 0.000 ;
  SIZE 88.240 BY 182.520 ;
  PIN vddio
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 7.000 171.090 76.510 172.520 ;
        RECT 7.000 79.905 8.430 171.090 ;
        RECT 14.300 165.925 48.885 167.285 ;
        RECT 14.300 156.525 15.660 165.925 ;
        RECT 47.525 156.525 48.885 165.925 ;
        RECT 14.300 155.165 48.885 156.525 ;
        RECT 15.005 106.480 51.690 121.685 ;
        RECT 15.005 103.880 67.505 106.480 ;
        RECT 15.005 97.510 67.505 100.110 ;
        RECT 15.570 93.640 50.130 97.510 ;
        RECT 15.570 84.605 50.130 88.765 ;
        RECT 75.080 79.905 76.510 171.090 ;
        RECT 7.000 78.475 76.510 79.905 ;
      LAYER li1 ;
        RECT 7.685 167.985 75.825 171.835 ;
        RECT 7.685 83.305 12.235 167.985 ;
        RECT 14.630 166.255 48.555 166.955 ;
        RECT 14.630 156.195 15.330 166.255 ;
        RECT 47.855 156.195 48.555 166.255 ;
        RECT 14.630 155.495 48.555 156.195 ;
        RECT 15.395 121.125 21.645 121.295 ;
        RECT 15.395 118.935 15.565 121.125 ;
        RECT 21.475 118.935 21.645 121.125 ;
        RECT 15.395 108.895 16.235 118.935 ;
        RECT 17.645 108.895 17.815 118.935 ;
        RECT 19.225 108.895 19.395 118.935 ;
        RECT 20.805 108.895 21.645 118.935 ;
        RECT 15.395 107.040 15.565 108.895 ;
        RECT 21.475 107.040 21.645 108.895 ;
        RECT 15.395 106.870 21.645 107.040 ;
        RECT 22.425 121.125 31.460 121.295 ;
        RECT 22.425 118.935 22.595 121.125 ;
        RECT 31.290 118.935 31.460 121.125 ;
        RECT 22.425 108.895 23.265 118.935 ;
        RECT 24.675 108.895 24.845 118.935 ;
        RECT 26.255 108.895 26.425 118.935 ;
        RECT 27.835 108.895 28.005 118.935 ;
        RECT 29.415 108.895 29.585 118.935 ;
        RECT 30.620 108.895 31.460 118.935 ;
        RECT 22.425 107.040 22.595 108.895 ;
        RECT 31.290 107.040 31.460 108.895 ;
        RECT 22.425 106.870 31.460 107.040 ;
        RECT 32.240 121.125 51.300 121.295 ;
        RECT 32.240 118.935 32.410 121.125 ;
        RECT 51.130 118.935 51.300 121.125 ;
        RECT 32.240 108.895 33.080 118.935 ;
        RECT 34.490 108.895 34.660 118.935 ;
        RECT 36.070 108.895 36.240 118.935 ;
        RECT 37.650 108.895 37.820 118.935 ;
        RECT 39.230 108.895 39.400 118.935 ;
        RECT 40.810 108.895 40.980 118.935 ;
        RECT 42.390 108.895 42.560 118.935 ;
        RECT 43.970 108.895 44.140 118.935 ;
        RECT 45.550 108.895 45.720 118.935 ;
        RECT 47.130 108.895 47.300 118.935 ;
        RECT 48.710 108.895 48.880 118.935 ;
        RECT 50.290 108.895 51.300 118.935 ;
        RECT 32.240 107.040 32.410 108.895 ;
        RECT 51.130 107.040 51.300 108.895 ;
        RECT 32.240 106.870 51.300 107.040 ;
        RECT 15.335 105.980 67.175 106.150 ;
        RECT 15.425 104.170 16.015 105.750 ;
        RECT 16.885 104.275 17.835 105.750 ;
        RECT 18.455 104.275 19.045 105.750 ;
        RECT 19.300 104.170 19.830 105.750 ;
        RECT 20.575 104.170 21.465 105.750 ;
        RECT 22.135 104.170 23.025 105.750 ;
        RECT 23.695 104.170 24.585 105.750 ;
        RECT 25.255 104.170 26.145 105.750 ;
        RECT 26.815 104.170 27.705 105.750 ;
        RECT 28.375 104.170 29.265 105.750 ;
        RECT 29.935 104.170 30.825 105.750 ;
        RECT 31.495 104.170 32.110 105.670 ;
        RECT 32.705 104.170 33.295 105.750 ;
        RECT 34.165 104.275 35.115 105.750 ;
        RECT 35.735 104.275 36.325 105.750 ;
        RECT 36.580 104.170 37.110 105.750 ;
        RECT 37.855 104.170 38.745 105.750 ;
        RECT 39.415 104.170 40.305 105.750 ;
        RECT 40.975 104.170 41.865 105.750 ;
        RECT 42.535 104.170 43.425 105.750 ;
        RECT 44.095 104.170 44.985 105.750 ;
        RECT 45.655 104.170 46.545 105.750 ;
        RECT 47.215 104.170 48.105 105.750 ;
        RECT 48.775 104.170 49.390 105.670 ;
        RECT 49.985 104.170 50.575 105.750 ;
        RECT 51.445 104.275 52.395 105.750 ;
        RECT 53.015 104.275 53.605 105.750 ;
        RECT 53.860 104.170 54.390 105.750 ;
        RECT 55.135 104.170 56.025 105.750 ;
        RECT 56.695 104.170 57.585 105.750 ;
        RECT 58.255 104.170 59.145 105.750 ;
        RECT 59.815 104.170 60.705 105.750 ;
        RECT 61.375 104.170 62.265 105.750 ;
        RECT 62.935 104.170 63.825 105.750 ;
        RECT 64.495 104.170 65.385 105.750 ;
        RECT 66.055 104.170 66.670 105.670 ;
        RECT 15.425 98.240 16.015 99.820 ;
        RECT 16.885 98.240 17.835 99.715 ;
        RECT 18.455 98.240 19.045 99.715 ;
        RECT 19.300 98.240 19.830 99.820 ;
        RECT 20.575 98.240 21.465 99.820 ;
        RECT 22.135 98.240 23.025 99.820 ;
        RECT 23.695 98.240 24.585 99.820 ;
        RECT 25.255 98.240 26.145 99.820 ;
        RECT 26.815 98.240 27.705 99.820 ;
        RECT 28.375 98.240 29.265 99.820 ;
        RECT 29.935 98.240 30.825 99.820 ;
        RECT 31.495 98.320 32.110 99.820 ;
        RECT 32.705 98.240 33.295 99.820 ;
        RECT 34.165 98.240 35.115 99.715 ;
        RECT 35.735 98.240 36.325 99.715 ;
        RECT 36.580 98.240 37.110 99.820 ;
        RECT 37.855 98.240 38.745 99.820 ;
        RECT 39.415 98.240 40.305 99.820 ;
        RECT 40.975 98.240 41.865 99.820 ;
        RECT 42.535 98.240 43.425 99.820 ;
        RECT 44.095 98.240 44.985 99.820 ;
        RECT 45.655 98.240 46.545 99.820 ;
        RECT 47.215 98.240 48.105 99.820 ;
        RECT 48.775 98.320 49.390 99.820 ;
        RECT 49.985 98.240 50.575 99.820 ;
        RECT 51.445 98.240 52.395 99.715 ;
        RECT 53.015 98.240 53.605 99.715 ;
        RECT 53.860 98.240 54.390 99.820 ;
        RECT 55.135 98.240 56.025 99.820 ;
        RECT 56.695 98.240 57.585 99.820 ;
        RECT 58.255 98.240 59.145 99.820 ;
        RECT 59.815 98.240 60.705 99.820 ;
        RECT 61.375 98.240 62.265 99.820 ;
        RECT 62.935 98.240 63.825 99.820 ;
        RECT 64.495 98.240 65.385 99.820 ;
        RECT 66.055 98.320 66.670 99.820 ;
        RECT 15.335 97.840 67.175 98.010 ;
        RECT 15.960 96.950 20.940 97.120 ;
        RECT 15.960 94.200 16.130 96.950 ;
        RECT 17.955 96.280 18.995 96.950 ;
        RECT 20.770 94.200 20.940 96.950 ;
        RECT 15.960 94.030 20.940 94.200 ;
        RECT 21.720 96.950 26.700 97.120 ;
        RECT 21.720 94.200 21.890 96.950 ;
        RECT 23.715 96.280 24.755 96.950 ;
        RECT 26.530 94.200 26.700 96.950 ;
        RECT 21.720 94.030 26.700 94.200 ;
        RECT 27.480 96.950 32.460 97.120 ;
        RECT 27.480 94.200 27.650 96.950 ;
        RECT 29.475 96.280 30.515 96.950 ;
        RECT 32.290 94.200 32.460 96.950 ;
        RECT 27.480 94.030 32.460 94.200 ;
        RECT 33.240 96.950 38.220 97.120 ;
        RECT 33.240 94.200 33.410 96.950 ;
        RECT 35.235 96.280 36.275 96.950 ;
        RECT 38.050 94.200 38.220 96.950 ;
        RECT 33.240 94.030 38.220 94.200 ;
        RECT 39.000 96.950 43.980 97.120 ;
        RECT 39.000 94.200 39.170 96.950 ;
        RECT 40.995 96.280 42.035 96.950 ;
        RECT 43.810 94.200 43.980 96.950 ;
        RECT 39.000 94.030 43.980 94.200 ;
        RECT 44.760 96.950 49.740 97.120 ;
        RECT 44.760 94.200 44.930 96.950 ;
        RECT 46.755 96.280 47.795 96.950 ;
        RECT 49.570 94.200 49.740 96.950 ;
        RECT 44.760 94.030 49.740 94.200 ;
        RECT 15.960 88.205 20.940 88.375 ;
        RECT 15.960 85.165 16.130 88.205 ;
        RECT 17.955 85.165 18.995 85.835 ;
        RECT 20.770 85.165 20.940 88.205 ;
        RECT 15.960 84.995 20.940 85.165 ;
        RECT 21.720 88.205 26.700 88.375 ;
        RECT 21.720 85.165 21.890 88.205 ;
        RECT 23.715 85.165 24.755 85.835 ;
        RECT 26.530 85.165 26.700 88.205 ;
        RECT 21.720 84.995 26.700 85.165 ;
        RECT 27.480 88.205 32.460 88.375 ;
        RECT 27.480 85.165 27.650 88.205 ;
        RECT 29.475 85.165 30.515 85.835 ;
        RECT 32.290 85.165 32.460 88.205 ;
        RECT 27.480 84.995 32.460 85.165 ;
        RECT 33.240 88.205 38.220 88.375 ;
        RECT 33.240 85.165 33.410 88.205 ;
        RECT 35.235 85.165 36.275 85.835 ;
        RECT 38.050 85.165 38.220 88.205 ;
        RECT 33.240 84.995 38.220 85.165 ;
        RECT 39.000 88.205 43.980 88.375 ;
        RECT 39.000 85.165 39.170 88.205 ;
        RECT 40.995 85.165 42.035 85.835 ;
        RECT 43.810 85.165 43.980 88.205 ;
        RECT 39.000 84.995 43.980 85.165 ;
        RECT 44.760 88.205 49.740 88.375 ;
        RECT 44.760 85.165 44.930 88.205 ;
        RECT 46.755 85.165 47.795 85.835 ;
        RECT 49.570 85.165 49.740 88.205 ;
        RECT 44.760 84.995 49.740 85.165 ;
        RECT 71.355 83.305 75.825 167.985 ;
        RECT 7.685 79.160 75.825 83.305 ;
      LAYER mcon ;
        RECT 15.830 166.545 16.000 166.715 ;
        RECT 16.190 166.545 16.360 166.715 ;
        RECT 16.550 166.545 16.720 166.715 ;
        RECT 16.910 166.545 17.080 166.715 ;
        RECT 17.270 166.545 17.440 166.715 ;
        RECT 17.630 166.545 17.800 166.715 ;
        RECT 17.990 166.545 18.160 166.715 ;
        RECT 18.350 166.545 18.520 166.715 ;
        RECT 18.710 166.545 18.880 166.715 ;
        RECT 19.070 166.545 19.240 166.715 ;
        RECT 19.430 166.545 19.600 166.715 ;
        RECT 19.790 166.545 19.960 166.715 ;
        RECT 20.315 166.545 20.485 166.715 ;
        RECT 20.675 166.545 20.845 166.715 ;
        RECT 21.035 166.545 21.205 166.715 ;
        RECT 21.395 166.545 21.565 166.715 ;
        RECT 21.755 166.545 21.925 166.715 ;
        RECT 22.115 166.545 22.285 166.715 ;
        RECT 22.475 166.545 22.645 166.715 ;
        RECT 22.835 166.545 23.005 166.715 ;
        RECT 23.195 166.545 23.365 166.715 ;
        RECT 23.555 166.545 23.725 166.715 ;
        RECT 23.915 166.545 24.085 166.715 ;
        RECT 24.275 166.545 24.445 166.715 ;
        RECT 24.780 166.545 24.950 166.715 ;
        RECT 25.140 166.545 25.310 166.715 ;
        RECT 25.500 166.545 25.670 166.715 ;
        RECT 25.860 166.545 26.030 166.715 ;
        RECT 26.220 166.545 26.390 166.715 ;
        RECT 26.580 166.545 26.750 166.715 ;
        RECT 26.940 166.545 27.110 166.715 ;
        RECT 27.300 166.545 27.470 166.715 ;
        RECT 27.660 166.545 27.830 166.715 ;
        RECT 28.020 166.545 28.190 166.715 ;
        RECT 28.380 166.545 28.550 166.715 ;
        RECT 28.740 166.545 28.910 166.715 ;
        RECT 29.265 166.545 29.435 166.715 ;
        RECT 29.625 166.545 29.795 166.715 ;
        RECT 29.985 166.545 30.155 166.715 ;
        RECT 30.345 166.545 30.515 166.715 ;
        RECT 30.705 166.545 30.875 166.715 ;
        RECT 31.065 166.545 31.235 166.715 ;
        RECT 31.425 166.545 31.595 166.715 ;
        RECT 31.785 166.545 31.955 166.715 ;
        RECT 32.555 166.545 32.725 166.715 ;
        RECT 32.915 166.545 33.085 166.715 ;
        RECT 33.275 166.545 33.445 166.715 ;
        RECT 33.635 166.545 33.805 166.715 ;
        RECT 33.995 166.545 34.165 166.715 ;
        RECT 34.355 166.545 34.525 166.715 ;
        RECT 34.715 166.545 34.885 166.715 ;
        RECT 35.075 166.545 35.245 166.715 ;
        RECT 35.435 166.545 35.605 166.715 ;
        RECT 35.795 166.545 35.965 166.715 ;
        RECT 36.155 166.545 36.325 166.715 ;
        RECT 36.515 166.545 36.685 166.715 ;
        RECT 37.040 166.545 37.210 166.715 ;
        RECT 37.400 166.545 37.570 166.715 ;
        RECT 37.760 166.545 37.930 166.715 ;
        RECT 38.120 166.545 38.290 166.715 ;
        RECT 38.480 166.545 38.650 166.715 ;
        RECT 38.840 166.545 39.010 166.715 ;
        RECT 39.200 166.545 39.370 166.715 ;
        RECT 39.560 166.545 39.730 166.715 ;
        RECT 39.920 166.545 40.090 166.715 ;
        RECT 40.280 166.545 40.450 166.715 ;
        RECT 40.640 166.545 40.810 166.715 ;
        RECT 41.000 166.545 41.170 166.715 ;
        RECT 41.505 166.545 41.675 166.715 ;
        RECT 41.865 166.545 42.035 166.715 ;
        RECT 42.225 166.545 42.395 166.715 ;
        RECT 42.585 166.545 42.755 166.715 ;
        RECT 42.945 166.545 43.115 166.715 ;
        RECT 43.305 166.545 43.475 166.715 ;
        RECT 43.665 166.545 43.835 166.715 ;
        RECT 44.025 166.545 44.195 166.715 ;
        RECT 44.385 166.545 44.555 166.715 ;
        RECT 44.745 166.545 44.915 166.715 ;
        RECT 45.105 166.545 45.275 166.715 ;
        RECT 45.465 166.545 45.635 166.715 ;
        RECT 45.990 166.545 46.160 166.715 ;
        RECT 46.350 166.545 46.520 166.715 ;
        RECT 46.710 166.545 46.880 166.715 ;
        RECT 47.070 166.545 47.240 166.715 ;
        RECT 47.430 166.545 47.600 166.715 ;
        RECT 14.895 165.170 15.065 165.340 ;
        RECT 14.895 164.810 15.065 164.980 ;
        RECT 14.895 164.450 15.065 164.620 ;
        RECT 14.895 164.090 15.065 164.260 ;
        RECT 14.895 163.730 15.065 163.900 ;
        RECT 14.895 163.370 15.065 163.540 ;
        RECT 14.895 163.010 15.065 163.180 ;
        RECT 14.895 162.650 15.065 162.820 ;
        RECT 14.895 162.290 15.065 162.460 ;
        RECT 14.895 161.930 15.065 162.100 ;
        RECT 14.895 161.570 15.065 161.740 ;
        RECT 14.895 161.210 15.065 161.380 ;
        RECT 14.895 160.850 15.065 161.020 ;
        RECT 14.895 160.490 15.065 160.660 ;
        RECT 14.895 160.130 15.065 160.300 ;
        RECT 14.895 159.770 15.065 159.940 ;
        RECT 14.895 159.410 15.065 159.580 ;
        RECT 14.895 159.050 15.065 159.220 ;
        RECT 14.895 158.690 15.065 158.860 ;
        RECT 14.895 158.330 15.065 158.500 ;
        RECT 14.895 157.970 15.065 158.140 ;
        RECT 14.895 157.610 15.065 157.780 ;
        RECT 14.895 157.250 15.065 157.420 ;
        RECT 14.895 156.890 15.065 157.060 ;
        RECT 14.895 156.530 15.065 156.700 ;
        RECT 48.100 165.170 48.270 165.340 ;
        RECT 48.100 164.810 48.270 164.980 ;
        RECT 48.100 164.450 48.270 164.620 ;
        RECT 48.100 164.090 48.270 164.260 ;
        RECT 48.100 163.730 48.270 163.900 ;
        RECT 48.100 163.370 48.270 163.540 ;
        RECT 48.100 163.010 48.270 163.180 ;
        RECT 48.100 162.650 48.270 162.820 ;
        RECT 48.100 162.290 48.270 162.460 ;
        RECT 48.100 161.930 48.270 162.100 ;
        RECT 48.100 161.570 48.270 161.740 ;
        RECT 48.100 161.210 48.270 161.380 ;
        RECT 48.100 160.850 48.270 161.020 ;
        RECT 48.100 160.490 48.270 160.660 ;
        RECT 48.100 160.130 48.270 160.300 ;
        RECT 48.100 159.770 48.270 159.940 ;
        RECT 48.100 159.410 48.270 159.580 ;
        RECT 48.100 159.050 48.270 159.220 ;
        RECT 48.100 158.690 48.270 158.860 ;
        RECT 48.100 158.330 48.270 158.500 ;
        RECT 48.100 157.970 48.270 158.140 ;
        RECT 48.100 157.610 48.270 157.780 ;
        RECT 48.100 157.250 48.270 157.420 ;
        RECT 48.100 156.890 48.270 157.060 ;
        RECT 48.100 156.530 48.270 156.700 ;
        RECT 15.830 155.755 16.000 155.925 ;
        RECT 16.190 155.755 16.360 155.925 ;
        RECT 16.550 155.755 16.720 155.925 ;
        RECT 16.910 155.755 17.080 155.925 ;
        RECT 17.270 155.755 17.440 155.925 ;
        RECT 17.630 155.755 17.800 155.925 ;
        RECT 17.990 155.755 18.160 155.925 ;
        RECT 18.350 155.755 18.520 155.925 ;
        RECT 18.710 155.755 18.880 155.925 ;
        RECT 19.070 155.755 19.240 155.925 ;
        RECT 19.430 155.755 19.600 155.925 ;
        RECT 19.790 155.755 19.960 155.925 ;
        RECT 20.315 155.755 20.485 155.925 ;
        RECT 20.675 155.755 20.845 155.925 ;
        RECT 21.035 155.755 21.205 155.925 ;
        RECT 21.395 155.755 21.565 155.925 ;
        RECT 21.755 155.755 21.925 155.925 ;
        RECT 22.115 155.755 22.285 155.925 ;
        RECT 22.475 155.755 22.645 155.925 ;
        RECT 22.835 155.755 23.005 155.925 ;
        RECT 23.195 155.755 23.365 155.925 ;
        RECT 23.555 155.755 23.725 155.925 ;
        RECT 23.915 155.755 24.085 155.925 ;
        RECT 24.275 155.755 24.445 155.925 ;
        RECT 24.780 155.755 24.950 155.925 ;
        RECT 25.140 155.755 25.310 155.925 ;
        RECT 25.500 155.755 25.670 155.925 ;
        RECT 25.860 155.755 26.030 155.925 ;
        RECT 26.220 155.755 26.390 155.925 ;
        RECT 26.580 155.755 26.750 155.925 ;
        RECT 26.940 155.755 27.110 155.925 ;
        RECT 27.300 155.755 27.470 155.925 ;
        RECT 27.660 155.755 27.830 155.925 ;
        RECT 28.020 155.755 28.190 155.925 ;
        RECT 28.380 155.755 28.550 155.925 ;
        RECT 28.740 155.755 28.910 155.925 ;
        RECT 29.265 155.755 29.435 155.925 ;
        RECT 29.625 155.755 29.795 155.925 ;
        RECT 29.985 155.755 30.155 155.925 ;
        RECT 30.345 155.755 30.515 155.925 ;
        RECT 30.705 155.755 30.875 155.925 ;
        RECT 31.065 155.755 31.235 155.925 ;
        RECT 31.425 155.755 31.595 155.925 ;
        RECT 31.785 155.755 31.955 155.925 ;
        RECT 32.325 155.755 32.495 155.925 ;
        RECT 32.685 155.755 32.855 155.925 ;
        RECT 33.045 155.755 33.215 155.925 ;
        RECT 33.405 155.755 33.575 155.925 ;
        RECT 33.765 155.755 33.935 155.925 ;
        RECT 34.125 155.755 34.295 155.925 ;
        RECT 34.485 155.755 34.655 155.925 ;
        RECT 34.845 155.755 35.015 155.925 ;
        RECT 35.205 155.755 35.375 155.925 ;
        RECT 35.565 155.755 35.735 155.925 ;
        RECT 35.925 155.755 36.095 155.925 ;
        RECT 36.285 155.755 36.455 155.925 ;
        RECT 36.810 155.755 36.980 155.925 ;
        RECT 37.170 155.755 37.340 155.925 ;
        RECT 37.530 155.755 37.700 155.925 ;
        RECT 37.890 155.755 38.060 155.925 ;
        RECT 38.250 155.755 38.420 155.925 ;
        RECT 38.610 155.755 38.780 155.925 ;
        RECT 38.970 155.755 39.140 155.925 ;
        RECT 39.330 155.755 39.500 155.925 ;
        RECT 39.690 155.755 39.860 155.925 ;
        RECT 40.050 155.755 40.220 155.925 ;
        RECT 40.410 155.755 40.580 155.925 ;
        RECT 40.770 155.755 40.940 155.925 ;
        RECT 41.275 155.755 41.445 155.925 ;
        RECT 41.635 155.755 41.805 155.925 ;
        RECT 41.995 155.755 42.165 155.925 ;
        RECT 42.355 155.755 42.525 155.925 ;
        RECT 42.715 155.755 42.885 155.925 ;
        RECT 43.075 155.755 43.245 155.925 ;
        RECT 43.435 155.755 43.605 155.925 ;
        RECT 43.795 155.755 43.965 155.925 ;
        RECT 44.155 155.755 44.325 155.925 ;
        RECT 44.515 155.755 44.685 155.925 ;
        RECT 44.875 155.755 45.045 155.925 ;
        RECT 45.235 155.755 45.405 155.925 ;
        RECT 45.760 155.755 45.930 155.925 ;
        RECT 46.120 155.755 46.290 155.925 ;
        RECT 46.480 155.755 46.650 155.925 ;
        RECT 46.840 155.755 47.010 155.925 ;
        RECT 47.200 155.755 47.370 155.925 ;
        RECT 9.625 130.080 9.795 130.250 ;
        RECT 9.985 130.080 10.155 130.250 ;
        RECT 10.345 130.080 10.515 130.250 ;
        RECT 10.705 130.080 10.875 130.250 ;
        RECT 11.065 130.080 11.235 130.250 ;
        RECT 11.425 130.080 11.595 130.250 ;
        RECT 9.625 129.565 9.795 129.735 ;
        RECT 9.985 129.565 10.155 129.735 ;
        RECT 10.345 129.565 10.515 129.735 ;
        RECT 10.705 129.565 10.875 129.735 ;
        RECT 11.065 129.565 11.235 129.735 ;
        RECT 11.425 129.565 11.595 129.735 ;
        RECT 9.625 129.110 9.795 129.280 ;
        RECT 9.985 129.110 10.155 129.280 ;
        RECT 10.345 129.110 10.515 129.280 ;
        RECT 10.705 129.110 10.875 129.280 ;
        RECT 11.065 129.110 11.235 129.280 ;
        RECT 11.425 129.110 11.595 129.280 ;
        RECT 9.625 128.595 9.795 128.765 ;
        RECT 9.985 128.595 10.155 128.765 ;
        RECT 10.345 128.595 10.515 128.765 ;
        RECT 10.705 128.595 10.875 128.765 ;
        RECT 11.065 128.595 11.235 128.765 ;
        RECT 11.425 128.595 11.595 128.765 ;
        RECT 9.625 128.085 9.795 128.255 ;
        RECT 9.985 128.085 10.155 128.255 ;
        RECT 10.345 128.085 10.515 128.255 ;
        RECT 10.705 128.085 10.875 128.255 ;
        RECT 11.065 128.085 11.235 128.255 ;
        RECT 11.425 128.085 11.595 128.255 ;
        RECT 9.625 127.565 9.795 127.735 ;
        RECT 9.985 127.565 10.155 127.735 ;
        RECT 10.345 127.565 10.515 127.735 ;
        RECT 10.705 127.565 10.875 127.735 ;
        RECT 11.065 127.565 11.235 127.735 ;
        RECT 11.425 127.565 11.595 127.735 ;
        RECT 9.625 127.115 9.795 127.285 ;
        RECT 9.985 127.115 10.155 127.285 ;
        RECT 10.345 127.115 10.515 127.285 ;
        RECT 10.705 127.115 10.875 127.285 ;
        RECT 11.065 127.115 11.235 127.285 ;
        RECT 11.425 127.115 11.595 127.285 ;
        RECT 9.625 126.600 9.795 126.770 ;
        RECT 9.985 126.600 10.155 126.770 ;
        RECT 10.345 126.600 10.515 126.770 ;
        RECT 10.705 126.600 10.875 126.770 ;
        RECT 11.065 126.600 11.235 126.770 ;
        RECT 11.425 126.600 11.595 126.770 ;
        RECT 9.625 126.125 9.795 126.295 ;
        RECT 9.985 126.125 10.155 126.295 ;
        RECT 10.345 126.125 10.515 126.295 ;
        RECT 10.705 126.125 10.875 126.295 ;
        RECT 11.065 126.125 11.235 126.295 ;
        RECT 11.425 126.125 11.595 126.295 ;
        RECT 9.625 125.605 9.795 125.775 ;
        RECT 9.985 125.605 10.155 125.775 ;
        RECT 10.345 125.605 10.515 125.775 ;
        RECT 10.705 125.605 10.875 125.775 ;
        RECT 11.065 125.605 11.235 125.775 ;
        RECT 11.425 125.605 11.595 125.775 ;
        RECT 72.665 130.245 72.835 130.415 ;
        RECT 73.025 130.245 73.195 130.415 ;
        RECT 73.385 130.245 73.555 130.415 ;
        RECT 73.745 130.245 73.915 130.415 ;
        RECT 74.105 130.245 74.275 130.415 ;
        RECT 74.465 130.245 74.635 130.415 ;
        RECT 72.665 129.730 72.835 129.900 ;
        RECT 73.025 129.730 73.195 129.900 ;
        RECT 73.385 129.730 73.555 129.900 ;
        RECT 73.745 129.730 73.915 129.900 ;
        RECT 74.105 129.730 74.275 129.900 ;
        RECT 74.465 129.730 74.635 129.900 ;
        RECT 72.665 129.275 72.835 129.445 ;
        RECT 73.025 129.275 73.195 129.445 ;
        RECT 73.385 129.275 73.555 129.445 ;
        RECT 73.745 129.275 73.915 129.445 ;
        RECT 74.105 129.275 74.275 129.445 ;
        RECT 74.465 129.275 74.635 129.445 ;
        RECT 72.665 128.760 72.835 128.930 ;
        RECT 73.025 128.760 73.195 128.930 ;
        RECT 73.385 128.760 73.555 128.930 ;
        RECT 73.745 128.760 73.915 128.930 ;
        RECT 74.105 128.760 74.275 128.930 ;
        RECT 74.465 128.760 74.635 128.930 ;
        RECT 72.665 128.250 72.835 128.420 ;
        RECT 73.025 128.250 73.195 128.420 ;
        RECT 73.385 128.250 73.555 128.420 ;
        RECT 73.745 128.250 73.915 128.420 ;
        RECT 74.105 128.250 74.275 128.420 ;
        RECT 74.465 128.250 74.635 128.420 ;
        RECT 72.665 127.730 72.835 127.900 ;
        RECT 73.025 127.730 73.195 127.900 ;
        RECT 73.385 127.730 73.555 127.900 ;
        RECT 73.745 127.730 73.915 127.900 ;
        RECT 74.105 127.730 74.275 127.900 ;
        RECT 74.465 127.730 74.635 127.900 ;
        RECT 72.665 127.280 72.835 127.450 ;
        RECT 73.025 127.280 73.195 127.450 ;
        RECT 73.385 127.280 73.555 127.450 ;
        RECT 73.745 127.280 73.915 127.450 ;
        RECT 74.105 127.280 74.275 127.450 ;
        RECT 74.465 127.280 74.635 127.450 ;
        RECT 72.665 126.765 72.835 126.935 ;
        RECT 73.025 126.765 73.195 126.935 ;
        RECT 73.385 126.765 73.555 126.935 ;
        RECT 73.745 126.765 73.915 126.935 ;
        RECT 74.105 126.765 74.275 126.935 ;
        RECT 74.465 126.765 74.635 126.935 ;
        RECT 72.665 126.290 72.835 126.460 ;
        RECT 73.025 126.290 73.195 126.460 ;
        RECT 73.385 126.290 73.555 126.460 ;
        RECT 73.745 126.290 73.915 126.460 ;
        RECT 74.105 126.290 74.275 126.460 ;
        RECT 74.465 126.290 74.635 126.460 ;
        RECT 72.665 125.770 72.835 125.940 ;
        RECT 73.025 125.770 73.195 125.940 ;
        RECT 73.385 125.770 73.555 125.940 ;
        RECT 73.745 125.770 73.915 125.940 ;
        RECT 74.105 125.770 74.275 125.940 ;
        RECT 74.465 125.770 74.635 125.940 ;
        RECT 15.660 118.510 15.830 118.680 ;
        RECT 16.065 118.510 16.235 118.680 ;
        RECT 15.660 118.150 15.830 118.320 ;
        RECT 16.065 118.150 16.235 118.320 ;
        RECT 15.660 117.790 15.830 117.960 ;
        RECT 16.065 117.790 16.235 117.960 ;
        RECT 15.660 114.465 15.830 114.635 ;
        RECT 16.065 114.410 16.235 114.580 ;
        RECT 15.660 114.105 15.830 114.275 ;
        RECT 16.065 114.050 16.235 114.220 ;
        RECT 16.065 113.690 16.235 113.860 ;
        RECT 15.660 110.740 15.830 110.910 ;
        RECT 16.065 110.615 16.235 110.785 ;
        RECT 15.660 110.380 15.830 110.550 ;
        RECT 16.065 110.255 16.235 110.425 ;
        RECT 15.660 110.020 15.830 110.190 ;
        RECT 16.065 109.895 16.235 110.065 ;
        RECT 17.645 118.510 17.815 118.680 ;
        RECT 17.645 118.150 17.815 118.320 ;
        RECT 17.645 117.790 17.815 117.960 ;
        RECT 17.645 114.410 17.815 114.580 ;
        RECT 17.645 114.050 17.815 114.220 ;
        RECT 17.645 113.690 17.815 113.860 ;
        RECT 17.645 110.615 17.815 110.785 ;
        RECT 17.645 110.255 17.815 110.425 ;
        RECT 17.645 109.895 17.815 110.065 ;
        RECT 19.225 118.510 19.395 118.680 ;
        RECT 19.225 118.150 19.395 118.320 ;
        RECT 19.225 117.790 19.395 117.960 ;
        RECT 19.225 114.410 19.395 114.580 ;
        RECT 19.225 114.050 19.395 114.220 ;
        RECT 19.225 113.690 19.395 113.860 ;
        RECT 19.225 110.615 19.395 110.785 ;
        RECT 19.225 110.255 19.395 110.425 ;
        RECT 19.225 109.895 19.395 110.065 ;
        RECT 20.805 118.510 20.975 118.680 ;
        RECT 21.180 118.510 21.350 118.680 ;
        RECT 20.805 118.150 20.975 118.320 ;
        RECT 21.180 118.150 21.350 118.320 ;
        RECT 20.805 117.790 20.975 117.960 ;
        RECT 21.180 117.790 21.350 117.960 ;
        RECT 20.805 114.410 20.975 114.580 ;
        RECT 21.180 114.465 21.350 114.635 ;
        RECT 20.805 114.050 20.975 114.220 ;
        RECT 21.180 114.105 21.350 114.275 ;
        RECT 20.805 113.690 20.975 113.860 ;
        RECT 20.805 110.615 20.975 110.785 ;
        RECT 21.180 110.740 21.350 110.910 ;
        RECT 20.805 110.255 20.975 110.425 ;
        RECT 21.180 110.380 21.350 110.550 ;
        RECT 20.805 109.895 20.975 110.065 ;
        RECT 21.180 110.020 21.350 110.190 ;
        RECT 22.690 118.510 22.860 118.680 ;
        RECT 23.095 118.510 23.265 118.680 ;
        RECT 22.690 118.150 22.860 118.320 ;
        RECT 23.095 118.150 23.265 118.320 ;
        RECT 22.690 117.790 22.860 117.960 ;
        RECT 23.095 117.790 23.265 117.960 ;
        RECT 22.690 114.500 22.860 114.670 ;
        RECT 23.095 114.410 23.265 114.580 ;
        RECT 22.690 114.140 22.860 114.310 ;
        RECT 23.095 114.050 23.265 114.220 ;
        RECT 22.690 113.780 22.860 113.950 ;
        RECT 23.095 113.690 23.265 113.860 ;
        RECT 22.690 110.690 22.860 110.860 ;
        RECT 23.095 110.615 23.265 110.785 ;
        RECT 22.690 110.330 22.860 110.500 ;
        RECT 23.095 110.255 23.265 110.425 ;
        RECT 22.690 109.970 22.860 110.140 ;
        RECT 23.095 109.895 23.265 110.065 ;
        RECT 24.675 118.510 24.845 118.680 ;
        RECT 24.675 118.150 24.845 118.320 ;
        RECT 24.675 117.790 24.845 117.960 ;
        RECT 24.675 114.410 24.845 114.580 ;
        RECT 24.675 114.050 24.845 114.220 ;
        RECT 24.675 113.690 24.845 113.860 ;
        RECT 24.675 110.615 24.845 110.785 ;
        RECT 24.675 110.255 24.845 110.425 ;
        RECT 24.675 109.895 24.845 110.065 ;
        RECT 26.255 118.510 26.425 118.680 ;
        RECT 26.255 118.150 26.425 118.320 ;
        RECT 26.255 117.790 26.425 117.960 ;
        RECT 26.255 114.410 26.425 114.580 ;
        RECT 26.255 114.050 26.425 114.220 ;
        RECT 26.255 113.690 26.425 113.860 ;
        RECT 26.255 110.615 26.425 110.785 ;
        RECT 26.255 110.255 26.425 110.425 ;
        RECT 26.255 109.895 26.425 110.065 ;
        RECT 27.835 118.510 28.005 118.680 ;
        RECT 27.835 118.150 28.005 118.320 ;
        RECT 27.835 117.790 28.005 117.960 ;
        RECT 27.835 114.410 28.005 114.580 ;
        RECT 27.835 114.050 28.005 114.220 ;
        RECT 27.835 113.690 28.005 113.860 ;
        RECT 27.835 110.615 28.005 110.785 ;
        RECT 27.835 110.255 28.005 110.425 ;
        RECT 27.835 109.895 28.005 110.065 ;
        RECT 29.415 118.510 29.585 118.680 ;
        RECT 29.415 118.150 29.585 118.320 ;
        RECT 29.415 117.790 29.585 117.960 ;
        RECT 29.415 114.410 29.585 114.580 ;
        RECT 29.415 114.050 29.585 114.220 ;
        RECT 29.415 113.690 29.585 113.860 ;
        RECT 29.415 110.615 29.585 110.785 ;
        RECT 29.415 110.255 29.585 110.425 ;
        RECT 29.415 109.895 29.585 110.065 ;
        RECT 30.995 118.510 31.165 118.680 ;
        RECT 30.995 118.150 31.165 118.320 ;
        RECT 30.995 117.790 31.165 117.960 ;
        RECT 30.995 114.500 31.165 114.670 ;
        RECT 30.995 114.140 31.165 114.310 ;
        RECT 30.995 113.780 31.165 113.950 ;
        RECT 30.995 110.740 31.165 110.910 ;
        RECT 30.995 110.380 31.165 110.550 ;
        RECT 30.995 110.020 31.165 110.190 ;
        RECT 32.505 118.510 32.675 118.680 ;
        RECT 32.910 118.510 33.080 118.680 ;
        RECT 32.505 118.150 32.675 118.320 ;
        RECT 32.910 118.150 33.080 118.320 ;
        RECT 32.505 117.790 32.675 117.960 ;
        RECT 32.910 117.790 33.080 117.960 ;
        RECT 32.505 114.480 32.675 114.650 ;
        RECT 32.910 114.410 33.080 114.580 ;
        RECT 32.505 114.120 32.675 114.290 ;
        RECT 32.910 114.050 33.080 114.220 ;
        RECT 32.505 113.760 32.675 113.930 ;
        RECT 32.910 113.690 33.080 113.860 ;
        RECT 32.505 110.740 32.675 110.910 ;
        RECT 32.910 110.615 33.080 110.785 ;
        RECT 32.505 110.380 32.675 110.550 ;
        RECT 32.910 110.255 33.080 110.425 ;
        RECT 32.505 110.020 32.675 110.190 ;
        RECT 32.910 109.895 33.080 110.065 ;
        RECT 34.490 118.510 34.660 118.680 ;
        RECT 34.490 118.150 34.660 118.320 ;
        RECT 34.490 117.790 34.660 117.960 ;
        RECT 34.490 114.410 34.660 114.580 ;
        RECT 34.490 114.050 34.660 114.220 ;
        RECT 34.490 113.690 34.660 113.860 ;
        RECT 34.490 110.615 34.660 110.785 ;
        RECT 34.490 110.255 34.660 110.425 ;
        RECT 34.490 109.895 34.660 110.065 ;
        RECT 36.070 118.510 36.240 118.680 ;
        RECT 36.070 118.150 36.240 118.320 ;
        RECT 36.070 117.790 36.240 117.960 ;
        RECT 36.070 114.410 36.240 114.580 ;
        RECT 36.070 114.050 36.240 114.220 ;
        RECT 36.070 113.690 36.240 113.860 ;
        RECT 36.070 110.615 36.240 110.785 ;
        RECT 36.070 110.255 36.240 110.425 ;
        RECT 36.070 109.895 36.240 110.065 ;
        RECT 37.650 118.510 37.820 118.680 ;
        RECT 37.650 118.150 37.820 118.320 ;
        RECT 37.650 117.790 37.820 117.960 ;
        RECT 37.650 114.410 37.820 114.580 ;
        RECT 37.650 114.050 37.820 114.220 ;
        RECT 37.650 113.690 37.820 113.860 ;
        RECT 37.650 110.615 37.820 110.785 ;
        RECT 37.650 110.255 37.820 110.425 ;
        RECT 37.650 109.895 37.820 110.065 ;
        RECT 39.230 118.510 39.400 118.680 ;
        RECT 39.230 118.150 39.400 118.320 ;
        RECT 39.230 117.790 39.400 117.960 ;
        RECT 39.230 114.410 39.400 114.580 ;
        RECT 39.230 114.050 39.400 114.220 ;
        RECT 39.230 113.690 39.400 113.860 ;
        RECT 39.230 110.615 39.400 110.785 ;
        RECT 39.230 110.255 39.400 110.425 ;
        RECT 39.230 109.895 39.400 110.065 ;
        RECT 40.810 118.510 40.980 118.680 ;
        RECT 40.810 118.150 40.980 118.320 ;
        RECT 40.810 117.790 40.980 117.960 ;
        RECT 40.810 114.410 40.980 114.580 ;
        RECT 40.810 114.050 40.980 114.220 ;
        RECT 40.810 113.690 40.980 113.860 ;
        RECT 40.810 110.615 40.980 110.785 ;
        RECT 40.810 110.255 40.980 110.425 ;
        RECT 40.810 109.895 40.980 110.065 ;
        RECT 42.390 118.510 42.560 118.680 ;
        RECT 42.390 118.150 42.560 118.320 ;
        RECT 42.390 117.790 42.560 117.960 ;
        RECT 42.390 114.410 42.560 114.580 ;
        RECT 42.390 114.050 42.560 114.220 ;
        RECT 42.390 113.690 42.560 113.860 ;
        RECT 42.390 110.615 42.560 110.785 ;
        RECT 42.390 110.255 42.560 110.425 ;
        RECT 42.390 109.895 42.560 110.065 ;
        RECT 43.970 118.510 44.140 118.680 ;
        RECT 43.970 118.150 44.140 118.320 ;
        RECT 43.970 117.790 44.140 117.960 ;
        RECT 43.970 114.410 44.140 114.580 ;
        RECT 43.970 114.050 44.140 114.220 ;
        RECT 43.970 113.690 44.140 113.860 ;
        RECT 43.970 110.615 44.140 110.785 ;
        RECT 43.970 110.255 44.140 110.425 ;
        RECT 43.970 109.895 44.140 110.065 ;
        RECT 45.550 118.510 45.720 118.680 ;
        RECT 45.550 118.150 45.720 118.320 ;
        RECT 45.550 117.790 45.720 117.960 ;
        RECT 45.550 114.410 45.720 114.580 ;
        RECT 45.550 114.050 45.720 114.220 ;
        RECT 45.550 113.690 45.720 113.860 ;
        RECT 45.550 110.615 45.720 110.785 ;
        RECT 45.550 110.255 45.720 110.425 ;
        RECT 45.550 109.895 45.720 110.065 ;
        RECT 47.130 118.510 47.300 118.680 ;
        RECT 47.130 118.150 47.300 118.320 ;
        RECT 47.130 117.790 47.300 117.960 ;
        RECT 47.130 114.410 47.300 114.580 ;
        RECT 47.130 114.050 47.300 114.220 ;
        RECT 47.130 113.690 47.300 113.860 ;
        RECT 47.130 110.615 47.300 110.785 ;
        RECT 47.130 110.255 47.300 110.425 ;
        RECT 47.130 109.895 47.300 110.065 ;
        RECT 48.710 118.510 48.880 118.680 ;
        RECT 48.710 118.150 48.880 118.320 ;
        RECT 48.710 117.790 48.880 117.960 ;
        RECT 48.710 114.410 48.880 114.580 ;
        RECT 48.710 114.050 48.880 114.220 ;
        RECT 48.710 113.690 48.880 113.860 ;
        RECT 48.710 110.615 48.880 110.785 ;
        RECT 48.710 110.255 48.880 110.425 ;
        RECT 48.710 109.895 48.880 110.065 ;
        RECT 50.290 118.510 50.460 118.680 ;
        RECT 50.835 118.510 51.005 118.680 ;
        RECT 50.290 118.150 50.460 118.320 ;
        RECT 50.835 118.150 51.005 118.320 ;
        RECT 50.290 117.790 50.460 117.960 ;
        RECT 50.835 117.790 51.005 117.960 ;
        RECT 50.290 114.410 50.460 114.580 ;
        RECT 50.835 114.435 51.005 114.605 ;
        RECT 50.290 114.050 50.460 114.220 ;
        RECT 50.835 114.075 51.005 114.245 ;
        RECT 50.290 113.690 50.460 113.860 ;
        RECT 50.835 113.715 51.005 113.885 ;
        RECT 50.290 110.615 50.460 110.785 ;
        RECT 50.835 110.740 51.005 110.910 ;
        RECT 50.290 110.255 50.460 110.425 ;
        RECT 50.835 110.380 51.005 110.550 ;
        RECT 50.290 109.895 50.460 110.065 ;
        RECT 50.835 110.020 51.005 110.190 ;
        RECT 15.490 105.980 15.660 106.150 ;
        RECT 15.970 105.980 16.140 106.150 ;
        RECT 16.450 105.980 16.620 106.150 ;
        RECT 16.930 105.980 17.100 106.150 ;
        RECT 17.410 105.980 17.580 106.150 ;
        RECT 17.890 105.980 18.060 106.150 ;
        RECT 18.370 105.980 18.540 106.150 ;
        RECT 18.850 105.980 19.020 106.150 ;
        RECT 19.330 105.980 19.500 106.150 ;
        RECT 19.810 105.980 19.980 106.150 ;
        RECT 20.290 105.980 20.460 106.150 ;
        RECT 20.770 105.980 20.940 106.150 ;
        RECT 21.250 105.980 21.420 106.150 ;
        RECT 21.730 105.980 21.900 106.150 ;
        RECT 22.210 105.980 22.380 106.150 ;
        RECT 22.690 105.980 22.860 106.150 ;
        RECT 23.170 105.980 23.340 106.150 ;
        RECT 23.650 105.980 23.820 106.150 ;
        RECT 24.130 105.980 24.300 106.150 ;
        RECT 24.610 105.980 24.780 106.150 ;
        RECT 25.090 105.980 25.260 106.150 ;
        RECT 25.570 105.980 25.740 106.150 ;
        RECT 26.050 105.980 26.220 106.150 ;
        RECT 26.530 105.980 26.700 106.150 ;
        RECT 27.010 105.980 27.180 106.150 ;
        RECT 27.490 105.980 27.660 106.150 ;
        RECT 27.970 105.980 28.140 106.150 ;
        RECT 28.450 105.980 28.620 106.150 ;
        RECT 28.930 105.980 29.100 106.150 ;
        RECT 29.410 105.980 29.580 106.150 ;
        RECT 29.890 105.980 30.060 106.150 ;
        RECT 30.370 105.980 30.540 106.150 ;
        RECT 30.850 105.980 31.020 106.150 ;
        RECT 31.330 105.980 31.500 106.150 ;
        RECT 31.810 105.980 31.980 106.150 ;
        RECT 32.290 105.980 32.460 106.150 ;
        RECT 32.770 105.980 32.940 106.150 ;
        RECT 33.250 105.980 33.420 106.150 ;
        RECT 33.730 105.980 33.900 106.150 ;
        RECT 34.210 105.980 34.380 106.150 ;
        RECT 34.690 105.980 34.860 106.150 ;
        RECT 35.170 105.980 35.340 106.150 ;
        RECT 35.650 105.980 35.820 106.150 ;
        RECT 36.130 105.980 36.300 106.150 ;
        RECT 36.610 105.980 36.780 106.150 ;
        RECT 37.090 105.980 37.260 106.150 ;
        RECT 37.570 105.980 37.740 106.150 ;
        RECT 38.050 105.980 38.220 106.150 ;
        RECT 38.530 105.980 38.700 106.150 ;
        RECT 39.010 105.980 39.180 106.150 ;
        RECT 39.490 105.980 39.660 106.150 ;
        RECT 39.970 105.980 40.140 106.150 ;
        RECT 40.450 105.980 40.620 106.150 ;
        RECT 40.930 105.980 41.100 106.150 ;
        RECT 41.410 105.980 41.580 106.150 ;
        RECT 41.890 105.980 42.060 106.150 ;
        RECT 42.370 105.980 42.540 106.150 ;
        RECT 42.850 105.980 43.020 106.150 ;
        RECT 43.330 105.980 43.500 106.150 ;
        RECT 43.810 105.980 43.980 106.150 ;
        RECT 44.290 105.980 44.460 106.150 ;
        RECT 44.770 105.980 44.940 106.150 ;
        RECT 45.250 105.980 45.420 106.150 ;
        RECT 45.730 105.980 45.900 106.150 ;
        RECT 46.210 105.980 46.380 106.150 ;
        RECT 46.690 105.980 46.860 106.150 ;
        RECT 47.170 105.980 47.340 106.150 ;
        RECT 47.650 105.980 47.820 106.150 ;
        RECT 48.130 105.980 48.300 106.150 ;
        RECT 48.610 105.980 48.780 106.150 ;
        RECT 49.090 105.980 49.260 106.150 ;
        RECT 49.570 105.980 49.740 106.150 ;
        RECT 50.050 105.980 50.220 106.150 ;
        RECT 50.530 105.980 50.700 106.150 ;
        RECT 51.010 105.980 51.180 106.150 ;
        RECT 51.490 105.980 51.660 106.150 ;
        RECT 51.970 105.980 52.140 106.150 ;
        RECT 52.450 105.980 52.620 106.150 ;
        RECT 52.930 105.980 53.100 106.150 ;
        RECT 53.410 105.980 53.580 106.150 ;
        RECT 53.890 105.980 54.060 106.150 ;
        RECT 54.370 105.980 54.540 106.150 ;
        RECT 54.850 105.980 55.020 106.150 ;
        RECT 55.330 105.980 55.500 106.150 ;
        RECT 55.810 105.980 55.980 106.150 ;
        RECT 56.290 105.980 56.460 106.150 ;
        RECT 56.770 105.980 56.940 106.150 ;
        RECT 57.250 105.980 57.420 106.150 ;
        RECT 57.730 105.980 57.900 106.150 ;
        RECT 58.210 105.980 58.380 106.150 ;
        RECT 58.690 105.980 58.860 106.150 ;
        RECT 59.170 105.980 59.340 106.150 ;
        RECT 59.650 105.980 59.820 106.150 ;
        RECT 60.130 105.980 60.300 106.150 ;
        RECT 60.610 105.980 60.780 106.150 ;
        RECT 61.090 105.980 61.260 106.150 ;
        RECT 61.570 105.980 61.740 106.150 ;
        RECT 62.050 105.980 62.220 106.150 ;
        RECT 62.530 105.980 62.700 106.150 ;
        RECT 63.010 105.980 63.180 106.150 ;
        RECT 63.490 105.980 63.660 106.150 ;
        RECT 63.970 105.980 64.140 106.150 ;
        RECT 64.450 105.980 64.620 106.150 ;
        RECT 64.930 105.980 65.100 106.150 ;
        RECT 65.410 105.980 65.580 106.150 ;
        RECT 65.890 105.980 66.060 106.150 ;
        RECT 66.370 105.980 66.540 106.150 ;
        RECT 66.850 105.980 67.020 106.150 ;
        RECT 15.455 105.500 15.625 105.670 ;
        RECT 15.815 105.500 15.985 105.670 ;
        RECT 16.915 105.500 17.085 105.670 ;
        RECT 17.275 105.500 17.445 105.670 ;
        RECT 17.635 105.500 17.805 105.670 ;
        RECT 18.485 105.500 18.655 105.670 ;
        RECT 18.845 105.500 19.015 105.670 ;
        RECT 19.300 105.470 19.470 105.640 ;
        RECT 19.660 105.470 19.830 105.640 ;
        RECT 20.575 105.470 20.745 105.640 ;
        RECT 20.935 105.470 21.105 105.640 ;
        RECT 21.295 105.470 21.465 105.640 ;
        RECT 22.135 105.470 22.305 105.640 ;
        RECT 22.495 105.470 22.665 105.640 ;
        RECT 22.855 105.470 23.025 105.640 ;
        RECT 23.695 105.470 23.865 105.640 ;
        RECT 24.055 105.470 24.225 105.640 ;
        RECT 24.415 105.470 24.585 105.640 ;
        RECT 25.255 105.470 25.425 105.640 ;
        RECT 25.615 105.470 25.785 105.640 ;
        RECT 25.975 105.470 26.145 105.640 ;
        RECT 26.815 105.470 26.985 105.640 ;
        RECT 27.175 105.470 27.345 105.640 ;
        RECT 27.535 105.470 27.705 105.640 ;
        RECT 28.375 105.470 28.545 105.640 ;
        RECT 28.735 105.470 28.905 105.640 ;
        RECT 29.095 105.470 29.265 105.640 ;
        RECT 29.935 105.470 30.105 105.640 ;
        RECT 30.295 105.470 30.465 105.640 ;
        RECT 30.655 105.470 30.825 105.640 ;
        RECT 31.540 105.470 31.710 105.640 ;
        RECT 31.900 105.470 32.070 105.640 ;
        RECT 32.735 105.500 32.905 105.670 ;
        RECT 33.095 105.500 33.265 105.670 ;
        RECT 34.195 105.500 34.365 105.670 ;
        RECT 34.555 105.500 34.725 105.670 ;
        RECT 34.915 105.500 35.085 105.670 ;
        RECT 35.765 105.500 35.935 105.670 ;
        RECT 36.125 105.500 36.295 105.670 ;
        RECT 36.580 105.470 36.750 105.640 ;
        RECT 36.940 105.470 37.110 105.640 ;
        RECT 37.855 105.470 38.025 105.640 ;
        RECT 38.215 105.470 38.385 105.640 ;
        RECT 38.575 105.470 38.745 105.640 ;
        RECT 39.415 105.470 39.585 105.640 ;
        RECT 39.775 105.470 39.945 105.640 ;
        RECT 40.135 105.470 40.305 105.640 ;
        RECT 40.975 105.470 41.145 105.640 ;
        RECT 41.335 105.470 41.505 105.640 ;
        RECT 41.695 105.470 41.865 105.640 ;
        RECT 42.535 105.470 42.705 105.640 ;
        RECT 42.895 105.470 43.065 105.640 ;
        RECT 43.255 105.470 43.425 105.640 ;
        RECT 44.095 105.470 44.265 105.640 ;
        RECT 44.455 105.470 44.625 105.640 ;
        RECT 44.815 105.470 44.985 105.640 ;
        RECT 45.655 105.470 45.825 105.640 ;
        RECT 46.015 105.470 46.185 105.640 ;
        RECT 46.375 105.470 46.545 105.640 ;
        RECT 47.215 105.470 47.385 105.640 ;
        RECT 47.575 105.470 47.745 105.640 ;
        RECT 47.935 105.470 48.105 105.640 ;
        RECT 48.820 105.470 48.990 105.640 ;
        RECT 49.180 105.470 49.350 105.640 ;
        RECT 50.015 105.500 50.185 105.670 ;
        RECT 50.375 105.500 50.545 105.670 ;
        RECT 51.475 105.500 51.645 105.670 ;
        RECT 51.835 105.500 52.005 105.670 ;
        RECT 52.195 105.500 52.365 105.670 ;
        RECT 53.045 105.500 53.215 105.670 ;
        RECT 53.405 105.500 53.575 105.670 ;
        RECT 53.860 105.470 54.030 105.640 ;
        RECT 54.220 105.470 54.390 105.640 ;
        RECT 55.135 105.470 55.305 105.640 ;
        RECT 55.495 105.470 55.665 105.640 ;
        RECT 55.855 105.470 56.025 105.640 ;
        RECT 56.695 105.470 56.865 105.640 ;
        RECT 57.055 105.470 57.225 105.640 ;
        RECT 57.415 105.470 57.585 105.640 ;
        RECT 58.255 105.470 58.425 105.640 ;
        RECT 58.615 105.470 58.785 105.640 ;
        RECT 58.975 105.470 59.145 105.640 ;
        RECT 59.815 105.470 59.985 105.640 ;
        RECT 60.175 105.470 60.345 105.640 ;
        RECT 60.535 105.470 60.705 105.640 ;
        RECT 61.375 105.470 61.545 105.640 ;
        RECT 61.735 105.470 61.905 105.640 ;
        RECT 62.095 105.470 62.265 105.640 ;
        RECT 62.935 105.470 63.105 105.640 ;
        RECT 63.295 105.470 63.465 105.640 ;
        RECT 63.655 105.470 63.825 105.640 ;
        RECT 64.495 105.470 64.665 105.640 ;
        RECT 64.855 105.470 65.025 105.640 ;
        RECT 65.215 105.470 65.385 105.640 ;
        RECT 66.100 105.470 66.270 105.640 ;
        RECT 66.460 105.470 66.630 105.640 ;
        RECT 15.455 98.320 15.625 98.490 ;
        RECT 15.815 98.320 15.985 98.490 ;
        RECT 16.915 98.320 17.085 98.490 ;
        RECT 17.275 98.320 17.445 98.490 ;
        RECT 17.635 98.320 17.805 98.490 ;
        RECT 18.485 98.320 18.655 98.490 ;
        RECT 18.845 98.320 19.015 98.490 ;
        RECT 19.300 98.350 19.470 98.520 ;
        RECT 19.660 98.350 19.830 98.520 ;
        RECT 20.575 98.350 20.745 98.520 ;
        RECT 20.935 98.350 21.105 98.520 ;
        RECT 21.295 98.350 21.465 98.520 ;
        RECT 22.135 98.350 22.305 98.520 ;
        RECT 22.495 98.350 22.665 98.520 ;
        RECT 22.855 98.350 23.025 98.520 ;
        RECT 23.695 98.350 23.865 98.520 ;
        RECT 24.055 98.350 24.225 98.520 ;
        RECT 24.415 98.350 24.585 98.520 ;
        RECT 25.255 98.350 25.425 98.520 ;
        RECT 25.615 98.350 25.785 98.520 ;
        RECT 25.975 98.350 26.145 98.520 ;
        RECT 26.815 98.350 26.985 98.520 ;
        RECT 27.175 98.350 27.345 98.520 ;
        RECT 27.535 98.350 27.705 98.520 ;
        RECT 28.375 98.350 28.545 98.520 ;
        RECT 28.735 98.350 28.905 98.520 ;
        RECT 29.095 98.350 29.265 98.520 ;
        RECT 29.935 98.350 30.105 98.520 ;
        RECT 30.295 98.350 30.465 98.520 ;
        RECT 30.655 98.350 30.825 98.520 ;
        RECT 31.540 98.350 31.710 98.520 ;
        RECT 31.900 98.350 32.070 98.520 ;
        RECT 32.735 98.320 32.905 98.490 ;
        RECT 33.095 98.320 33.265 98.490 ;
        RECT 34.195 98.320 34.365 98.490 ;
        RECT 34.555 98.320 34.725 98.490 ;
        RECT 34.915 98.320 35.085 98.490 ;
        RECT 35.765 98.320 35.935 98.490 ;
        RECT 36.125 98.320 36.295 98.490 ;
        RECT 36.580 98.350 36.750 98.520 ;
        RECT 36.940 98.350 37.110 98.520 ;
        RECT 37.855 98.350 38.025 98.520 ;
        RECT 38.215 98.350 38.385 98.520 ;
        RECT 38.575 98.350 38.745 98.520 ;
        RECT 39.415 98.350 39.585 98.520 ;
        RECT 39.775 98.350 39.945 98.520 ;
        RECT 40.135 98.350 40.305 98.520 ;
        RECT 40.975 98.350 41.145 98.520 ;
        RECT 41.335 98.350 41.505 98.520 ;
        RECT 41.695 98.350 41.865 98.520 ;
        RECT 42.535 98.350 42.705 98.520 ;
        RECT 42.895 98.350 43.065 98.520 ;
        RECT 43.255 98.350 43.425 98.520 ;
        RECT 44.095 98.350 44.265 98.520 ;
        RECT 44.455 98.350 44.625 98.520 ;
        RECT 44.815 98.350 44.985 98.520 ;
        RECT 45.655 98.350 45.825 98.520 ;
        RECT 46.015 98.350 46.185 98.520 ;
        RECT 46.375 98.350 46.545 98.520 ;
        RECT 47.215 98.350 47.385 98.520 ;
        RECT 47.575 98.350 47.745 98.520 ;
        RECT 47.935 98.350 48.105 98.520 ;
        RECT 48.820 98.350 48.990 98.520 ;
        RECT 49.180 98.350 49.350 98.520 ;
        RECT 50.015 98.320 50.185 98.490 ;
        RECT 50.375 98.320 50.545 98.490 ;
        RECT 51.475 98.320 51.645 98.490 ;
        RECT 51.835 98.320 52.005 98.490 ;
        RECT 52.195 98.320 52.365 98.490 ;
        RECT 53.045 98.320 53.215 98.490 ;
        RECT 53.405 98.320 53.575 98.490 ;
        RECT 53.860 98.350 54.030 98.520 ;
        RECT 54.220 98.350 54.390 98.520 ;
        RECT 55.135 98.350 55.305 98.520 ;
        RECT 55.495 98.350 55.665 98.520 ;
        RECT 55.855 98.350 56.025 98.520 ;
        RECT 56.695 98.350 56.865 98.520 ;
        RECT 57.055 98.350 57.225 98.520 ;
        RECT 57.415 98.350 57.585 98.520 ;
        RECT 58.255 98.350 58.425 98.520 ;
        RECT 58.615 98.350 58.785 98.520 ;
        RECT 58.975 98.350 59.145 98.520 ;
        RECT 59.815 98.350 59.985 98.520 ;
        RECT 60.175 98.350 60.345 98.520 ;
        RECT 60.535 98.350 60.705 98.520 ;
        RECT 61.375 98.350 61.545 98.520 ;
        RECT 61.735 98.350 61.905 98.520 ;
        RECT 62.095 98.350 62.265 98.520 ;
        RECT 62.935 98.350 63.105 98.520 ;
        RECT 63.295 98.350 63.465 98.520 ;
        RECT 63.655 98.350 63.825 98.520 ;
        RECT 64.495 98.350 64.665 98.520 ;
        RECT 64.855 98.350 65.025 98.520 ;
        RECT 65.215 98.350 65.385 98.520 ;
        RECT 66.100 98.350 66.270 98.520 ;
        RECT 66.460 98.350 66.630 98.520 ;
        RECT 15.490 97.840 15.660 98.010 ;
        RECT 15.970 97.840 16.140 98.010 ;
        RECT 16.450 97.840 16.620 98.010 ;
        RECT 16.930 97.840 17.100 98.010 ;
        RECT 17.410 97.840 17.580 98.010 ;
        RECT 17.890 97.840 18.060 98.010 ;
        RECT 18.370 97.840 18.540 98.010 ;
        RECT 18.850 97.840 19.020 98.010 ;
        RECT 19.330 97.840 19.500 98.010 ;
        RECT 19.810 97.840 19.980 98.010 ;
        RECT 20.290 97.840 20.460 98.010 ;
        RECT 20.770 97.840 20.940 98.010 ;
        RECT 21.250 97.840 21.420 98.010 ;
        RECT 21.730 97.840 21.900 98.010 ;
        RECT 22.210 97.840 22.380 98.010 ;
        RECT 22.690 97.840 22.860 98.010 ;
        RECT 23.170 97.840 23.340 98.010 ;
        RECT 23.650 97.840 23.820 98.010 ;
        RECT 24.130 97.840 24.300 98.010 ;
        RECT 24.610 97.840 24.780 98.010 ;
        RECT 25.090 97.840 25.260 98.010 ;
        RECT 25.570 97.840 25.740 98.010 ;
        RECT 26.050 97.840 26.220 98.010 ;
        RECT 26.530 97.840 26.700 98.010 ;
        RECT 27.010 97.840 27.180 98.010 ;
        RECT 27.490 97.840 27.660 98.010 ;
        RECT 27.970 97.840 28.140 98.010 ;
        RECT 28.450 97.840 28.620 98.010 ;
        RECT 28.930 97.840 29.100 98.010 ;
        RECT 29.410 97.840 29.580 98.010 ;
        RECT 29.890 97.840 30.060 98.010 ;
        RECT 30.370 97.840 30.540 98.010 ;
        RECT 30.850 97.840 31.020 98.010 ;
        RECT 31.330 97.840 31.500 98.010 ;
        RECT 31.810 97.840 31.980 98.010 ;
        RECT 32.290 97.840 32.460 98.010 ;
        RECT 32.770 97.840 32.940 98.010 ;
        RECT 33.250 97.840 33.420 98.010 ;
        RECT 33.730 97.840 33.900 98.010 ;
        RECT 34.210 97.840 34.380 98.010 ;
        RECT 34.690 97.840 34.860 98.010 ;
        RECT 35.170 97.840 35.340 98.010 ;
        RECT 35.650 97.840 35.820 98.010 ;
        RECT 36.130 97.840 36.300 98.010 ;
        RECT 36.610 97.840 36.780 98.010 ;
        RECT 37.090 97.840 37.260 98.010 ;
        RECT 37.570 97.840 37.740 98.010 ;
        RECT 38.050 97.840 38.220 98.010 ;
        RECT 38.530 97.840 38.700 98.010 ;
        RECT 39.010 97.840 39.180 98.010 ;
        RECT 39.490 97.840 39.660 98.010 ;
        RECT 39.970 97.840 40.140 98.010 ;
        RECT 40.450 97.840 40.620 98.010 ;
        RECT 40.930 97.840 41.100 98.010 ;
        RECT 41.410 97.840 41.580 98.010 ;
        RECT 41.890 97.840 42.060 98.010 ;
        RECT 42.370 97.840 42.540 98.010 ;
        RECT 42.850 97.840 43.020 98.010 ;
        RECT 43.330 97.840 43.500 98.010 ;
        RECT 43.810 97.840 43.980 98.010 ;
        RECT 44.290 97.840 44.460 98.010 ;
        RECT 44.770 97.840 44.940 98.010 ;
        RECT 45.250 97.840 45.420 98.010 ;
        RECT 45.730 97.840 45.900 98.010 ;
        RECT 46.210 97.840 46.380 98.010 ;
        RECT 46.690 97.840 46.860 98.010 ;
        RECT 47.170 97.840 47.340 98.010 ;
        RECT 47.650 97.840 47.820 98.010 ;
        RECT 48.130 97.840 48.300 98.010 ;
        RECT 48.610 97.840 48.780 98.010 ;
        RECT 49.090 97.840 49.260 98.010 ;
        RECT 49.570 97.840 49.740 98.010 ;
        RECT 50.050 97.840 50.220 98.010 ;
        RECT 50.530 97.840 50.700 98.010 ;
        RECT 51.010 97.840 51.180 98.010 ;
        RECT 51.490 97.840 51.660 98.010 ;
        RECT 51.970 97.840 52.140 98.010 ;
        RECT 52.450 97.840 52.620 98.010 ;
        RECT 52.930 97.840 53.100 98.010 ;
        RECT 53.410 97.840 53.580 98.010 ;
        RECT 53.890 97.840 54.060 98.010 ;
        RECT 54.370 97.840 54.540 98.010 ;
        RECT 54.850 97.840 55.020 98.010 ;
        RECT 55.330 97.840 55.500 98.010 ;
        RECT 55.810 97.840 55.980 98.010 ;
        RECT 56.290 97.840 56.460 98.010 ;
        RECT 56.770 97.840 56.940 98.010 ;
        RECT 57.250 97.840 57.420 98.010 ;
        RECT 57.730 97.840 57.900 98.010 ;
        RECT 58.210 97.840 58.380 98.010 ;
        RECT 58.690 97.840 58.860 98.010 ;
        RECT 59.170 97.840 59.340 98.010 ;
        RECT 59.650 97.840 59.820 98.010 ;
        RECT 60.130 97.840 60.300 98.010 ;
        RECT 60.610 97.840 60.780 98.010 ;
        RECT 61.090 97.840 61.260 98.010 ;
        RECT 61.570 97.840 61.740 98.010 ;
        RECT 62.050 97.840 62.220 98.010 ;
        RECT 62.530 97.840 62.700 98.010 ;
        RECT 63.010 97.840 63.180 98.010 ;
        RECT 63.490 97.840 63.660 98.010 ;
        RECT 63.970 97.840 64.140 98.010 ;
        RECT 64.450 97.840 64.620 98.010 ;
        RECT 64.930 97.840 65.100 98.010 ;
        RECT 65.410 97.840 65.580 98.010 ;
        RECT 65.890 97.840 66.060 98.010 ;
        RECT 66.370 97.840 66.540 98.010 ;
        RECT 66.850 97.840 67.020 98.010 ;
        RECT 18.190 96.950 18.360 97.120 ;
        RECT 18.550 96.950 18.720 97.120 ;
        RECT 18.190 96.280 18.360 96.450 ;
        RECT 18.550 96.280 18.720 96.450 ;
        RECT 23.950 96.950 24.120 97.120 ;
        RECT 24.310 96.950 24.480 97.120 ;
        RECT 23.950 96.280 24.120 96.450 ;
        RECT 24.310 96.280 24.480 96.450 ;
        RECT 29.710 96.950 29.880 97.120 ;
        RECT 30.070 96.950 30.240 97.120 ;
        RECT 29.710 96.280 29.880 96.450 ;
        RECT 30.070 96.280 30.240 96.450 ;
        RECT 35.470 96.950 35.640 97.120 ;
        RECT 35.830 96.950 36.000 97.120 ;
        RECT 35.470 96.280 35.640 96.450 ;
        RECT 35.830 96.280 36.000 96.450 ;
        RECT 41.230 96.950 41.400 97.120 ;
        RECT 41.590 96.950 41.760 97.120 ;
        RECT 41.230 96.280 41.400 96.450 ;
        RECT 41.590 96.280 41.760 96.450 ;
        RECT 46.990 96.950 47.160 97.120 ;
        RECT 47.350 96.950 47.520 97.120 ;
        RECT 46.990 96.280 47.160 96.450 ;
        RECT 47.350 96.280 47.520 96.450 ;
        RECT 18.330 85.395 18.500 85.565 ;
        RECT 18.690 85.395 18.860 85.565 ;
        RECT 18.330 84.995 18.500 85.165 ;
        RECT 18.690 84.995 18.860 85.165 ;
        RECT 24.090 85.395 24.260 85.565 ;
        RECT 24.450 85.395 24.620 85.565 ;
        RECT 24.090 84.995 24.260 85.165 ;
        RECT 24.450 84.995 24.620 85.165 ;
        RECT 29.850 85.395 30.020 85.565 ;
        RECT 30.210 85.395 30.380 85.565 ;
        RECT 29.850 84.995 30.020 85.165 ;
        RECT 30.210 84.995 30.380 85.165 ;
        RECT 35.610 85.395 35.780 85.565 ;
        RECT 35.970 85.395 36.140 85.565 ;
        RECT 35.610 84.995 35.780 85.165 ;
        RECT 35.970 84.995 36.140 85.165 ;
        RECT 41.370 85.395 41.540 85.565 ;
        RECT 41.730 85.395 41.900 85.565 ;
        RECT 41.370 84.995 41.540 85.165 ;
        RECT 41.730 84.995 41.900 85.165 ;
        RECT 47.130 85.395 47.300 85.565 ;
        RECT 47.490 85.395 47.660 85.565 ;
        RECT 47.130 84.995 47.300 85.165 ;
        RECT 47.490 84.995 47.660 85.165 ;
      LAYER met1 ;
        RECT 14.630 166.255 48.550 166.955 ;
        RECT 14.630 156.195 15.330 166.255 ;
        RECT 47.850 156.195 48.550 166.255 ;
        RECT 14.630 155.960 48.550 156.195 ;
        RECT 0.000 123.160 88.240 155.960 ;
        RECT 11.175 117.685 51.310 118.915 ;
        RECT 11.175 113.585 51.310 114.815 ;
        RECT 11.175 109.790 51.310 111.020 ;
        RECT 13.815 105.440 74.810 106.180 ;
        RECT 14.110 96.805 75.150 98.550 ;
        RECT 17.975 96.200 18.975 96.805 ;
        RECT 23.735 96.200 24.735 96.805 ;
        RECT 29.495 96.200 30.495 96.805 ;
        RECT 35.255 96.200 36.255 96.805 ;
        RECT 41.015 96.200 42.015 96.805 ;
        RECT 46.775 96.200 47.775 96.805 ;
        RECT 17.975 85.160 18.975 85.795 ;
        RECT 23.735 85.160 24.735 85.795 ;
        RECT 29.495 85.160 30.495 85.795 ;
        RECT 35.255 85.160 36.255 85.795 ;
        RECT 41.015 85.160 42.015 85.795 ;
        RECT 46.775 85.160 47.775 85.795 ;
        RECT 17.005 83.910 75.345 85.160 ;
      LAYER via ;
        RECT 70.940 132.385 71.200 132.645 ;
        RECT 71.280 132.385 71.540 132.645 ;
        RECT 71.600 132.385 71.860 132.645 ;
        RECT 72.005 132.385 72.265 132.645 ;
        RECT 72.345 132.385 72.605 132.645 ;
        RECT 72.665 132.385 72.925 132.645 ;
        RECT 73.150 132.385 73.410 132.645 ;
        RECT 73.490 132.385 73.750 132.645 ;
        RECT 73.810 132.385 74.070 132.645 ;
        RECT 74.215 132.385 74.475 132.645 ;
        RECT 74.555 132.385 74.815 132.645 ;
        RECT 70.940 132.060 71.200 132.320 ;
        RECT 71.280 132.060 71.540 132.320 ;
        RECT 71.600 132.060 71.860 132.320 ;
        RECT 72.005 132.060 72.265 132.320 ;
        RECT 72.345 132.060 72.605 132.320 ;
        RECT 72.665 132.060 72.925 132.320 ;
        RECT 73.150 132.060 73.410 132.320 ;
        RECT 73.490 132.060 73.750 132.320 ;
        RECT 73.810 132.060 74.070 132.320 ;
        RECT 74.215 132.060 74.475 132.320 ;
        RECT 74.555 132.060 74.815 132.320 ;
        RECT 70.940 131.730 71.200 131.990 ;
        RECT 71.280 131.730 71.540 131.990 ;
        RECT 71.600 131.730 71.860 131.990 ;
        RECT 72.005 131.730 72.265 131.990 ;
        RECT 72.345 131.730 72.605 131.990 ;
        RECT 72.665 131.730 72.925 131.990 ;
        RECT 73.150 131.730 73.410 131.990 ;
        RECT 73.490 131.730 73.750 131.990 ;
        RECT 73.810 131.730 74.070 131.990 ;
        RECT 74.215 131.730 74.475 131.990 ;
        RECT 74.555 131.730 74.815 131.990 ;
        RECT 70.940 131.330 71.200 131.590 ;
        RECT 71.280 131.330 71.540 131.590 ;
        RECT 71.600 131.330 71.860 131.590 ;
        RECT 72.005 131.330 72.265 131.590 ;
        RECT 72.345 131.330 72.605 131.590 ;
        RECT 72.665 131.330 72.925 131.590 ;
        RECT 73.150 131.330 73.410 131.590 ;
        RECT 73.490 131.330 73.750 131.590 ;
        RECT 73.810 131.330 74.070 131.590 ;
        RECT 74.215 131.330 74.475 131.590 ;
        RECT 74.555 131.330 74.815 131.590 ;
        RECT 70.940 131.005 71.200 131.265 ;
        RECT 71.280 131.005 71.540 131.265 ;
        RECT 71.600 131.005 71.860 131.265 ;
        RECT 72.005 131.005 72.265 131.265 ;
        RECT 72.345 131.005 72.605 131.265 ;
        RECT 72.665 131.005 72.925 131.265 ;
        RECT 73.150 131.005 73.410 131.265 ;
        RECT 73.490 131.005 73.750 131.265 ;
        RECT 73.810 131.005 74.070 131.265 ;
        RECT 74.215 131.005 74.475 131.265 ;
        RECT 74.555 131.005 74.815 131.265 ;
        RECT 70.940 130.675 71.200 130.935 ;
        RECT 71.280 130.675 71.540 130.935 ;
        RECT 71.600 130.675 71.860 130.935 ;
        RECT 72.005 130.675 72.265 130.935 ;
        RECT 72.345 130.675 72.605 130.935 ;
        RECT 72.665 130.675 72.925 130.935 ;
        RECT 73.150 130.675 73.410 130.935 ;
        RECT 73.490 130.675 73.750 130.935 ;
        RECT 73.810 130.675 74.070 130.935 ;
        RECT 74.215 130.675 74.475 130.935 ;
        RECT 74.555 130.675 74.815 130.935 ;
        RECT 70.940 130.205 71.200 130.465 ;
        RECT 71.280 130.205 71.540 130.465 ;
        RECT 71.600 130.205 71.860 130.465 ;
        RECT 72.005 130.205 72.265 130.465 ;
        RECT 72.345 130.205 72.605 130.465 ;
        RECT 72.665 130.205 72.925 130.465 ;
        RECT 73.150 130.205 73.410 130.465 ;
        RECT 73.490 130.205 73.750 130.465 ;
        RECT 73.810 130.205 74.070 130.465 ;
        RECT 74.215 130.205 74.475 130.465 ;
        RECT 74.555 130.205 74.815 130.465 ;
        RECT 70.940 129.880 71.200 130.140 ;
        RECT 71.280 129.880 71.540 130.140 ;
        RECT 71.600 129.880 71.860 130.140 ;
        RECT 72.005 129.880 72.265 130.140 ;
        RECT 72.345 129.880 72.605 130.140 ;
        RECT 72.665 129.880 72.925 130.140 ;
        RECT 73.150 129.880 73.410 130.140 ;
        RECT 73.490 129.880 73.750 130.140 ;
        RECT 73.810 129.880 74.070 130.140 ;
        RECT 74.215 129.880 74.475 130.140 ;
        RECT 74.555 129.880 74.815 130.140 ;
        RECT 70.940 129.550 71.200 129.810 ;
        RECT 71.280 129.550 71.540 129.810 ;
        RECT 71.600 129.550 71.860 129.810 ;
        RECT 72.005 129.550 72.265 129.810 ;
        RECT 72.345 129.550 72.605 129.810 ;
        RECT 72.665 129.550 72.925 129.810 ;
        RECT 73.150 129.550 73.410 129.810 ;
        RECT 73.490 129.550 73.750 129.810 ;
        RECT 73.810 129.550 74.070 129.810 ;
        RECT 74.215 129.550 74.475 129.810 ;
        RECT 74.555 129.550 74.815 129.810 ;
        RECT 70.940 129.150 71.200 129.410 ;
        RECT 71.280 129.150 71.540 129.410 ;
        RECT 71.600 129.150 71.860 129.410 ;
        RECT 72.005 129.150 72.265 129.410 ;
        RECT 72.345 129.150 72.605 129.410 ;
        RECT 72.665 129.150 72.925 129.410 ;
        RECT 73.150 129.150 73.410 129.410 ;
        RECT 73.490 129.150 73.750 129.410 ;
        RECT 73.810 129.150 74.070 129.410 ;
        RECT 74.215 129.150 74.475 129.410 ;
        RECT 74.555 129.150 74.815 129.410 ;
        RECT 70.940 128.825 71.200 129.085 ;
        RECT 71.280 128.825 71.540 129.085 ;
        RECT 71.600 128.825 71.860 129.085 ;
        RECT 72.005 128.825 72.265 129.085 ;
        RECT 72.345 128.825 72.605 129.085 ;
        RECT 72.665 128.825 72.925 129.085 ;
        RECT 73.150 128.825 73.410 129.085 ;
        RECT 73.490 128.825 73.750 129.085 ;
        RECT 73.810 128.825 74.070 129.085 ;
        RECT 74.215 128.825 74.475 129.085 ;
        RECT 74.555 128.825 74.815 129.085 ;
        RECT 70.940 128.495 71.200 128.755 ;
        RECT 71.280 128.495 71.540 128.755 ;
        RECT 71.600 128.495 71.860 128.755 ;
        RECT 72.005 128.495 72.265 128.755 ;
        RECT 72.345 128.495 72.605 128.755 ;
        RECT 72.665 128.495 72.925 128.755 ;
        RECT 73.150 128.495 73.410 128.755 ;
        RECT 73.490 128.495 73.750 128.755 ;
        RECT 73.810 128.495 74.070 128.755 ;
        RECT 74.215 128.495 74.475 128.755 ;
        RECT 74.555 128.495 74.815 128.755 ;
        RECT 70.940 127.965 71.200 128.225 ;
        RECT 71.280 127.965 71.540 128.225 ;
        RECT 71.600 127.965 71.860 128.225 ;
        RECT 72.005 127.965 72.265 128.225 ;
        RECT 72.345 127.965 72.605 128.225 ;
        RECT 72.665 127.965 72.925 128.225 ;
        RECT 73.150 127.965 73.410 128.225 ;
        RECT 73.490 127.965 73.750 128.225 ;
        RECT 73.810 127.965 74.070 128.225 ;
        RECT 74.215 127.965 74.475 128.225 ;
        RECT 74.555 127.965 74.815 128.225 ;
        RECT 13.555 127.690 13.815 127.950 ;
        RECT 13.895 127.690 14.155 127.950 ;
        RECT 14.215 127.690 14.475 127.950 ;
        RECT 70.940 127.640 71.200 127.900 ;
        RECT 71.280 127.640 71.540 127.900 ;
        RECT 71.600 127.640 71.860 127.900 ;
        RECT 72.005 127.640 72.265 127.900 ;
        RECT 72.345 127.640 72.605 127.900 ;
        RECT 72.665 127.640 72.925 127.900 ;
        RECT 73.150 127.640 73.410 127.900 ;
        RECT 73.490 127.640 73.750 127.900 ;
        RECT 73.810 127.640 74.070 127.900 ;
        RECT 74.215 127.640 74.475 127.900 ;
        RECT 74.555 127.640 74.815 127.900 ;
        RECT 13.555 127.365 13.815 127.625 ;
        RECT 13.895 127.365 14.155 127.625 ;
        RECT 14.215 127.365 14.475 127.625 ;
        RECT 70.940 127.310 71.200 127.570 ;
        RECT 71.280 127.310 71.540 127.570 ;
        RECT 71.600 127.310 71.860 127.570 ;
        RECT 72.005 127.310 72.265 127.570 ;
        RECT 72.345 127.310 72.605 127.570 ;
        RECT 72.665 127.310 72.925 127.570 ;
        RECT 73.150 127.310 73.410 127.570 ;
        RECT 73.490 127.310 73.750 127.570 ;
        RECT 73.810 127.310 74.070 127.570 ;
        RECT 74.215 127.310 74.475 127.570 ;
        RECT 74.555 127.310 74.815 127.570 ;
        RECT 13.555 127.035 13.815 127.295 ;
        RECT 13.895 127.035 14.155 127.295 ;
        RECT 14.215 127.035 14.475 127.295 ;
        RECT 70.940 126.910 71.200 127.170 ;
        RECT 71.280 126.910 71.540 127.170 ;
        RECT 71.600 126.910 71.860 127.170 ;
        RECT 72.005 126.910 72.265 127.170 ;
        RECT 72.345 126.910 72.605 127.170 ;
        RECT 72.665 126.910 72.925 127.170 ;
        RECT 73.150 126.910 73.410 127.170 ;
        RECT 73.490 126.910 73.750 127.170 ;
        RECT 73.810 126.910 74.070 127.170 ;
        RECT 74.215 126.910 74.475 127.170 ;
        RECT 74.555 126.910 74.815 127.170 ;
        RECT 13.555 126.635 13.815 126.895 ;
        RECT 13.895 126.635 14.155 126.895 ;
        RECT 14.215 126.635 14.475 126.895 ;
        RECT 70.940 126.585 71.200 126.845 ;
        RECT 71.280 126.585 71.540 126.845 ;
        RECT 71.600 126.585 71.860 126.845 ;
        RECT 72.005 126.585 72.265 126.845 ;
        RECT 72.345 126.585 72.605 126.845 ;
        RECT 72.665 126.585 72.925 126.845 ;
        RECT 73.150 126.585 73.410 126.845 ;
        RECT 73.490 126.585 73.750 126.845 ;
        RECT 73.810 126.585 74.070 126.845 ;
        RECT 74.215 126.585 74.475 126.845 ;
        RECT 74.555 126.585 74.815 126.845 ;
        RECT 13.555 126.310 13.815 126.570 ;
        RECT 13.895 126.310 14.155 126.570 ;
        RECT 14.215 126.310 14.475 126.570 ;
        RECT 70.940 126.255 71.200 126.515 ;
        RECT 71.280 126.255 71.540 126.515 ;
        RECT 71.600 126.255 71.860 126.515 ;
        RECT 72.005 126.255 72.265 126.515 ;
        RECT 72.345 126.255 72.605 126.515 ;
        RECT 72.665 126.255 72.925 126.515 ;
        RECT 73.150 126.255 73.410 126.515 ;
        RECT 73.490 126.255 73.750 126.515 ;
        RECT 73.810 126.255 74.070 126.515 ;
        RECT 74.215 126.255 74.475 126.515 ;
        RECT 74.555 126.255 74.815 126.515 ;
        RECT 13.555 125.980 13.815 126.240 ;
        RECT 13.895 125.980 14.155 126.240 ;
        RECT 14.215 125.980 14.475 126.240 ;
        RECT 70.940 125.785 71.200 126.045 ;
        RECT 71.280 125.785 71.540 126.045 ;
        RECT 71.600 125.785 71.860 126.045 ;
        RECT 72.005 125.785 72.265 126.045 ;
        RECT 72.345 125.785 72.605 126.045 ;
        RECT 72.665 125.785 72.925 126.045 ;
        RECT 73.150 125.785 73.410 126.045 ;
        RECT 73.490 125.785 73.750 126.045 ;
        RECT 73.810 125.785 74.070 126.045 ;
        RECT 74.215 125.785 74.475 126.045 ;
        RECT 74.555 125.785 74.815 126.045 ;
        RECT 13.555 125.510 13.815 125.770 ;
        RECT 13.895 125.510 14.155 125.770 ;
        RECT 14.215 125.510 14.475 125.770 ;
        RECT 70.940 125.460 71.200 125.720 ;
        RECT 71.280 125.460 71.540 125.720 ;
        RECT 71.600 125.460 71.860 125.720 ;
        RECT 72.005 125.460 72.265 125.720 ;
        RECT 72.345 125.460 72.605 125.720 ;
        RECT 72.665 125.460 72.925 125.720 ;
        RECT 73.150 125.460 73.410 125.720 ;
        RECT 73.490 125.460 73.750 125.720 ;
        RECT 73.810 125.460 74.070 125.720 ;
        RECT 74.215 125.460 74.475 125.720 ;
        RECT 74.555 125.460 74.815 125.720 ;
        RECT 13.555 125.185 13.815 125.445 ;
        RECT 13.895 125.185 14.155 125.445 ;
        RECT 14.215 125.185 14.475 125.445 ;
        RECT 70.940 125.130 71.200 125.390 ;
        RECT 71.280 125.130 71.540 125.390 ;
        RECT 71.600 125.130 71.860 125.390 ;
        RECT 72.005 125.130 72.265 125.390 ;
        RECT 72.345 125.130 72.605 125.390 ;
        RECT 72.665 125.130 72.925 125.390 ;
        RECT 73.150 125.130 73.410 125.390 ;
        RECT 73.490 125.130 73.750 125.390 ;
        RECT 73.810 125.130 74.070 125.390 ;
        RECT 74.215 125.130 74.475 125.390 ;
        RECT 74.555 125.130 74.815 125.390 ;
        RECT 13.555 124.855 13.815 125.115 ;
        RECT 13.895 124.855 14.155 125.115 ;
        RECT 14.215 124.855 14.475 125.115 ;
        RECT 70.940 124.730 71.200 124.990 ;
        RECT 71.280 124.730 71.540 124.990 ;
        RECT 71.600 124.730 71.860 124.990 ;
        RECT 72.005 124.730 72.265 124.990 ;
        RECT 72.345 124.730 72.605 124.990 ;
        RECT 72.665 124.730 72.925 124.990 ;
        RECT 73.150 124.730 73.410 124.990 ;
        RECT 73.490 124.730 73.750 124.990 ;
        RECT 73.810 124.730 74.070 124.990 ;
        RECT 74.215 124.730 74.475 124.990 ;
        RECT 74.555 124.730 74.815 124.990 ;
        RECT 13.555 124.455 13.815 124.715 ;
        RECT 13.895 124.455 14.155 124.715 ;
        RECT 14.215 124.455 14.475 124.715 ;
        RECT 70.940 124.405 71.200 124.665 ;
        RECT 71.280 124.405 71.540 124.665 ;
        RECT 71.600 124.405 71.860 124.665 ;
        RECT 72.005 124.405 72.265 124.665 ;
        RECT 72.345 124.405 72.605 124.665 ;
        RECT 72.665 124.405 72.925 124.665 ;
        RECT 73.150 124.405 73.410 124.665 ;
        RECT 73.490 124.405 73.750 124.665 ;
        RECT 73.810 124.405 74.070 124.665 ;
        RECT 74.215 124.405 74.475 124.665 ;
        RECT 74.555 124.405 74.815 124.665 ;
        RECT 13.555 124.130 13.815 124.390 ;
        RECT 13.895 124.130 14.155 124.390 ;
        RECT 14.215 124.130 14.475 124.390 ;
        RECT 70.940 124.075 71.200 124.335 ;
        RECT 71.280 124.075 71.540 124.335 ;
        RECT 71.600 124.075 71.860 124.335 ;
        RECT 72.005 124.075 72.265 124.335 ;
        RECT 72.345 124.075 72.605 124.335 ;
        RECT 72.665 124.075 72.925 124.335 ;
        RECT 73.150 124.075 73.410 124.335 ;
        RECT 73.490 124.075 73.750 124.335 ;
        RECT 73.810 124.075 74.070 124.335 ;
        RECT 74.215 124.075 74.475 124.335 ;
        RECT 74.555 124.075 74.815 124.335 ;
        RECT 13.555 123.800 13.815 124.060 ;
        RECT 13.895 123.800 14.155 124.060 ;
        RECT 14.215 123.800 14.475 124.060 ;
        RECT 13.265 118.485 13.525 118.745 ;
        RECT 13.605 118.485 13.865 118.745 ;
        RECT 13.925 118.485 14.185 118.745 ;
        RECT 14.330 118.485 14.590 118.745 ;
        RECT 14.670 118.485 14.930 118.745 ;
        RECT 13.265 118.160 13.525 118.420 ;
        RECT 13.605 118.160 13.865 118.420 ;
        RECT 13.925 118.160 14.185 118.420 ;
        RECT 14.330 118.160 14.590 118.420 ;
        RECT 14.670 118.160 14.930 118.420 ;
        RECT 13.265 117.830 13.525 118.090 ;
        RECT 13.605 117.830 13.865 118.090 ;
        RECT 13.925 117.830 14.185 118.090 ;
        RECT 14.330 117.830 14.590 118.090 ;
        RECT 14.670 117.830 14.930 118.090 ;
        RECT 13.265 114.420 13.525 114.680 ;
        RECT 13.605 114.420 13.865 114.680 ;
        RECT 13.925 114.420 14.185 114.680 ;
        RECT 14.330 114.420 14.590 114.680 ;
        RECT 14.670 114.420 14.930 114.680 ;
        RECT 13.265 114.095 13.525 114.355 ;
        RECT 13.605 114.095 13.865 114.355 ;
        RECT 13.925 114.095 14.185 114.355 ;
        RECT 14.330 114.095 14.590 114.355 ;
        RECT 14.670 114.095 14.930 114.355 ;
        RECT 13.265 113.765 13.525 114.025 ;
        RECT 13.605 113.765 13.865 114.025 ;
        RECT 13.925 113.765 14.185 114.025 ;
        RECT 14.330 113.765 14.590 114.025 ;
        RECT 14.670 113.765 14.930 114.025 ;
        RECT 13.265 110.555 13.525 110.815 ;
        RECT 13.605 110.555 13.865 110.815 ;
        RECT 13.925 110.555 14.185 110.815 ;
        RECT 14.330 110.555 14.590 110.815 ;
        RECT 14.670 110.555 14.930 110.815 ;
        RECT 13.265 110.230 13.525 110.490 ;
        RECT 13.605 110.230 13.865 110.490 ;
        RECT 13.925 110.230 14.185 110.490 ;
        RECT 14.330 110.230 14.590 110.490 ;
        RECT 14.670 110.230 14.930 110.490 ;
        RECT 13.265 109.900 13.525 110.160 ;
        RECT 13.605 109.900 13.865 110.160 ;
        RECT 13.925 109.900 14.185 110.160 ;
        RECT 14.330 109.900 14.590 110.160 ;
        RECT 14.670 109.900 14.930 110.160 ;
        RECT 71.015 105.815 71.275 106.075 ;
        RECT 71.355 105.815 71.615 106.075 ;
        RECT 71.675 105.815 71.935 106.075 ;
        RECT 72.080 105.815 72.340 106.075 ;
        RECT 72.420 105.815 72.680 106.075 ;
        RECT 72.740 105.815 73.000 106.075 ;
        RECT 73.210 105.815 73.470 106.075 ;
        RECT 73.550 105.815 73.810 106.075 ;
        RECT 73.870 105.815 74.130 106.075 ;
        RECT 74.275 105.815 74.535 106.075 ;
        RECT 71.015 105.490 71.275 105.750 ;
        RECT 71.355 105.490 71.615 105.750 ;
        RECT 71.675 105.490 71.935 105.750 ;
        RECT 72.080 105.490 72.340 105.750 ;
        RECT 72.420 105.490 72.680 105.750 ;
        RECT 72.740 105.490 73.000 105.750 ;
        RECT 73.210 105.490 73.470 105.750 ;
        RECT 73.550 105.490 73.810 105.750 ;
        RECT 73.870 105.490 74.130 105.750 ;
        RECT 74.275 105.490 74.535 105.750 ;
        RECT 71.015 97.850 71.275 98.110 ;
        RECT 71.355 97.850 71.615 98.110 ;
        RECT 71.675 97.850 71.935 98.110 ;
        RECT 72.080 97.850 72.340 98.110 ;
        RECT 72.420 97.850 72.680 98.110 ;
        RECT 72.740 97.850 73.000 98.110 ;
        RECT 73.210 97.850 73.470 98.110 ;
        RECT 73.550 97.850 73.810 98.110 ;
        RECT 73.870 97.850 74.130 98.110 ;
        RECT 74.275 97.850 74.535 98.110 ;
        RECT 71.015 97.525 71.275 97.785 ;
        RECT 71.355 97.525 71.615 97.785 ;
        RECT 71.675 97.525 71.935 97.785 ;
        RECT 72.080 97.525 72.340 97.785 ;
        RECT 72.420 97.525 72.680 97.785 ;
        RECT 72.740 97.525 73.000 97.785 ;
        RECT 73.210 97.525 73.470 97.785 ;
        RECT 73.550 97.525 73.810 97.785 ;
        RECT 73.870 97.525 74.130 97.785 ;
        RECT 74.275 97.525 74.535 97.785 ;
        RECT 71.015 97.195 71.275 97.455 ;
        RECT 71.355 97.195 71.615 97.455 ;
        RECT 71.675 97.195 71.935 97.455 ;
        RECT 72.080 97.195 72.340 97.455 ;
        RECT 72.420 97.195 72.680 97.455 ;
        RECT 72.740 97.195 73.000 97.455 ;
        RECT 73.210 97.195 73.470 97.455 ;
        RECT 73.550 97.195 73.810 97.455 ;
        RECT 73.870 97.195 74.130 97.455 ;
        RECT 74.275 97.195 74.535 97.455 ;
        RECT 71.015 84.740 71.275 85.000 ;
        RECT 71.355 84.740 71.615 85.000 ;
        RECT 71.675 84.740 71.935 85.000 ;
        RECT 72.080 84.740 72.340 85.000 ;
        RECT 72.420 84.740 72.680 85.000 ;
        RECT 72.740 84.740 73.000 85.000 ;
        RECT 73.210 84.740 73.470 85.000 ;
        RECT 73.550 84.740 73.810 85.000 ;
        RECT 73.870 84.740 74.130 85.000 ;
        RECT 74.275 84.740 74.535 85.000 ;
        RECT 71.015 84.415 71.275 84.675 ;
        RECT 71.355 84.415 71.615 84.675 ;
        RECT 71.675 84.415 71.935 84.675 ;
        RECT 72.080 84.415 72.340 84.675 ;
        RECT 72.420 84.415 72.680 84.675 ;
        RECT 72.740 84.415 73.000 84.675 ;
        RECT 73.210 84.415 73.470 84.675 ;
        RECT 73.550 84.415 73.810 84.675 ;
        RECT 73.870 84.415 74.130 84.675 ;
        RECT 74.275 84.415 74.535 84.675 ;
        RECT 71.015 84.085 71.275 84.345 ;
        RECT 71.355 84.085 71.615 84.345 ;
        RECT 71.675 84.085 71.935 84.345 ;
        RECT 72.080 84.085 72.340 84.345 ;
        RECT 72.420 84.085 72.680 84.345 ;
        RECT 72.740 84.085 73.000 84.345 ;
        RECT 73.210 84.085 73.470 84.345 ;
        RECT 73.550 84.085 73.810 84.345 ;
        RECT 73.870 84.085 74.130 84.345 ;
        RECT 74.275 84.085 74.535 84.345 ;
      LAYER met2 ;
        RECT 13.040 109.285 15.040 151.575 ;
        RECT 70.725 82.635 75.080 156.530 ;
    END
  END vddio
  PIN vssio
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 16.070 156.970 47.080 165.480 ;
        RECT 53.790 119.030 60.420 119.580 ;
        RECT 53.790 117.105 54.340 119.030 ;
        RECT 59.870 117.105 60.420 119.030 ;
        RECT 53.790 112.345 60.420 117.105 ;
        RECT 53.790 110.405 54.340 112.345 ;
        RECT 59.870 110.405 60.420 112.345 ;
        RECT 53.790 109.855 60.420 110.405 ;
        RECT 61.720 119.030 70.720 119.580 ;
        RECT 61.720 117.105 62.270 119.030 ;
        RECT 70.170 117.105 70.720 119.030 ;
        RECT 61.720 112.345 70.720 117.105 ;
        RECT 61.720 110.405 62.270 112.345 ;
        RECT 70.170 110.405 70.720 112.345 ;
        RECT 61.720 109.855 70.720 110.405 ;
        RECT 15.485 102.210 19.155 103.410 ;
        RECT 19.205 102.210 32.200 103.580 ;
        RECT 32.765 102.210 36.435 103.410 ;
        RECT 36.485 102.210 49.480 103.580 ;
        RECT 50.045 102.210 53.715 103.410 ;
        RECT 53.765 102.210 66.760 103.580 ;
        RECT 15.205 101.780 67.305 102.210 ;
        RECT 15.485 100.580 19.155 101.780 ;
        RECT 19.205 100.410 32.200 101.780 ;
        RECT 32.765 100.580 36.435 101.780 ;
        RECT 36.485 100.410 49.480 101.780 ;
        RECT 50.045 100.580 53.715 101.780 ;
        RECT 53.765 100.410 66.760 101.780 ;
        RECT 51.715 94.940 70.195 95.490 ;
        RECT 15.750 92.760 21.120 93.310 ;
        RECT 15.750 89.965 16.300 92.760 ;
        RECT 17.785 89.965 19.045 92.760 ;
        RECT 20.570 89.965 21.120 92.760 ;
        RECT 15.750 89.415 21.120 89.965 ;
        RECT 21.510 92.760 26.880 93.310 ;
        RECT 21.510 89.965 22.060 92.760 ;
        RECT 23.545 89.965 24.805 92.760 ;
        RECT 26.330 89.965 26.880 92.760 ;
        RECT 21.510 89.415 26.880 89.965 ;
        RECT 27.270 92.760 32.640 93.310 ;
        RECT 27.270 89.965 27.820 92.760 ;
        RECT 29.305 89.965 30.565 92.760 ;
        RECT 32.090 89.965 32.640 92.760 ;
        RECT 27.270 89.415 32.640 89.965 ;
        RECT 33.030 92.760 38.400 93.310 ;
        RECT 33.030 89.965 33.580 92.760 ;
        RECT 35.065 89.965 36.325 92.760 ;
        RECT 37.850 89.965 38.400 92.760 ;
        RECT 33.030 89.415 38.400 89.965 ;
        RECT 38.790 92.760 44.160 93.310 ;
        RECT 38.790 89.965 39.340 92.760 ;
        RECT 40.825 89.965 42.085 92.760 ;
        RECT 43.610 89.965 44.160 92.760 ;
        RECT 38.790 89.415 44.160 89.965 ;
        RECT 44.550 92.760 49.920 93.310 ;
        RECT 44.550 89.965 45.100 92.760 ;
        RECT 46.585 89.965 47.845 92.760 ;
        RECT 49.370 89.965 49.920 92.760 ;
        RECT 44.550 89.415 49.920 89.965 ;
        RECT 51.715 93.000 52.265 94.940 ;
        RECT 69.645 93.000 70.195 94.940 ;
        RECT 51.715 88.240 70.195 93.000 ;
        RECT 51.715 86.315 52.265 88.240 ;
        RECT 69.645 86.315 70.195 88.240 ;
        RECT 51.715 85.765 70.195 86.315 ;
      LAYER li1 ;
        RECT 16.240 164.155 31.265 165.310 ;
        RECT 16.240 158.315 17.960 164.155 ;
        RECT 21.030 158.315 22.020 164.155 ;
        RECT 25.060 158.315 26.050 164.155 ;
        RECT 29.030 158.315 31.265 164.155 ;
        RECT 16.240 158.150 31.265 158.315 ;
        RECT 31.885 164.155 46.910 165.310 ;
        RECT 31.885 158.315 34.120 164.155 ;
        RECT 37.100 158.315 38.090 164.155 ;
        RECT 41.130 158.315 42.120 164.155 ;
        RECT 45.190 158.315 46.910 164.155 ;
        RECT 31.885 158.150 46.910 158.315 ;
        RECT 16.240 157.140 31.250 158.150 ;
        RECT 31.900 157.140 46.910 158.150 ;
        RECT 53.980 119.220 60.230 119.390 ;
        RECT 53.980 116.995 54.150 119.220 ;
        RECT 60.060 116.995 60.230 119.220 ;
        RECT 53.980 112.455 54.820 116.995 ;
        RECT 56.230 112.455 56.400 116.995 ;
        RECT 57.810 112.455 57.980 116.995 ;
        RECT 59.390 112.455 60.230 116.995 ;
        RECT 53.980 110.215 54.150 112.455 ;
        RECT 60.060 110.215 60.230 112.455 ;
        RECT 53.980 110.045 60.230 110.215 ;
        RECT 61.910 119.220 70.530 119.390 ;
        RECT 61.910 116.995 62.080 119.220 ;
        RECT 61.910 112.455 62.750 116.995 ;
        RECT 64.160 112.455 64.330 116.995 ;
        RECT 65.740 112.455 65.910 116.995 ;
        RECT 67.320 112.455 67.490 116.995 ;
        RECT 68.900 112.455 69.070 116.995 ;
        RECT 61.910 110.215 62.080 112.455 ;
        RECT 70.360 110.215 70.530 119.220 ;
        RECT 61.910 110.045 70.530 110.215 ;
        RECT 15.425 102.360 16.015 103.320 ;
        RECT 16.805 102.360 17.755 103.045 ;
        RECT 18.715 102.360 19.045 103.320 ;
        RECT 19.270 102.370 19.805 103.470 ;
        RECT 20.575 102.370 21.465 103.390 ;
        RECT 22.135 102.370 23.025 103.390 ;
        RECT 23.695 102.370 24.585 103.390 ;
        RECT 25.255 102.370 26.145 103.390 ;
        RECT 26.815 102.370 27.705 103.390 ;
        RECT 28.375 102.370 29.265 103.390 ;
        RECT 29.935 102.370 30.825 103.390 ;
        RECT 31.495 102.370 32.110 103.390 ;
        RECT 32.705 102.360 33.295 103.320 ;
        RECT 34.085 102.360 35.035 103.045 ;
        RECT 35.995 102.360 36.325 103.320 ;
        RECT 36.550 102.370 37.085 103.470 ;
        RECT 37.855 102.370 38.745 103.390 ;
        RECT 39.415 102.370 40.305 103.390 ;
        RECT 40.975 102.370 41.865 103.390 ;
        RECT 42.535 102.370 43.425 103.390 ;
        RECT 44.095 102.370 44.985 103.390 ;
        RECT 45.655 102.370 46.545 103.390 ;
        RECT 47.215 102.370 48.105 103.390 ;
        RECT 48.775 102.370 49.390 103.390 ;
        RECT 49.985 102.360 50.575 103.320 ;
        RECT 51.365 102.360 52.315 103.045 ;
        RECT 53.275 102.360 53.605 103.320 ;
        RECT 53.830 102.370 54.365 103.470 ;
        RECT 55.135 102.370 56.025 103.390 ;
        RECT 56.695 102.370 57.585 103.390 ;
        RECT 58.255 102.370 59.145 103.390 ;
        RECT 59.815 102.370 60.705 103.390 ;
        RECT 61.375 102.370 62.265 103.390 ;
        RECT 62.935 102.370 63.825 103.390 ;
        RECT 64.495 102.370 65.385 103.390 ;
        RECT 66.055 102.370 66.670 103.390 ;
        RECT 15.335 101.910 67.175 102.080 ;
        RECT 15.425 100.670 16.015 101.630 ;
        RECT 16.805 100.945 17.755 101.630 ;
        RECT 18.715 100.670 19.045 101.630 ;
        RECT 19.270 100.520 19.805 101.620 ;
        RECT 20.575 100.600 21.465 101.620 ;
        RECT 22.135 100.600 23.025 101.620 ;
        RECT 23.695 100.600 24.585 101.620 ;
        RECT 25.255 100.600 26.145 101.620 ;
        RECT 26.815 100.600 27.705 101.620 ;
        RECT 28.375 100.600 29.265 101.620 ;
        RECT 29.935 100.600 30.825 101.620 ;
        RECT 31.495 100.600 32.110 101.620 ;
        RECT 32.705 100.670 33.295 101.630 ;
        RECT 34.085 100.945 35.035 101.630 ;
        RECT 35.995 100.670 36.325 101.630 ;
        RECT 36.550 100.520 37.085 101.620 ;
        RECT 37.855 100.600 38.745 101.620 ;
        RECT 39.415 100.600 40.305 101.620 ;
        RECT 40.975 100.600 41.865 101.620 ;
        RECT 42.535 100.600 43.425 101.620 ;
        RECT 44.095 100.600 44.985 101.620 ;
        RECT 45.655 100.600 46.545 101.620 ;
        RECT 47.215 100.600 48.105 101.620 ;
        RECT 48.775 100.600 49.390 101.620 ;
        RECT 49.985 100.670 50.575 101.630 ;
        RECT 51.365 100.945 52.315 101.630 ;
        RECT 53.275 100.670 53.605 101.630 ;
        RECT 53.830 100.520 54.365 101.620 ;
        RECT 55.135 100.600 56.025 101.620 ;
        RECT 56.695 100.600 57.585 101.620 ;
        RECT 58.255 100.600 59.145 101.620 ;
        RECT 59.815 100.600 60.705 101.620 ;
        RECT 61.375 100.600 62.265 101.620 ;
        RECT 62.935 100.600 63.825 101.620 ;
        RECT 64.495 100.600 65.385 101.620 ;
        RECT 66.055 100.600 66.670 101.620 ;
        RECT 51.905 95.130 70.005 95.300 ;
        RECT 15.770 92.950 21.100 93.120 ;
        RECT 15.770 91.385 16.110 92.950 ;
        RECT 17.895 91.385 18.935 91.525 ;
        RECT 20.760 91.385 21.100 92.950 ;
        RECT 15.770 91.215 21.100 91.385 ;
        RECT 15.770 89.775 16.110 91.215 ;
        RECT 17.895 91.065 18.935 91.215 ;
        RECT 20.760 89.775 21.100 91.215 ;
        RECT 15.770 89.605 21.100 89.775 ;
        RECT 21.530 92.950 26.860 93.120 ;
        RECT 21.530 91.385 21.870 92.950 ;
        RECT 23.655 91.385 24.695 91.525 ;
        RECT 26.520 91.385 26.860 92.950 ;
        RECT 21.530 91.215 26.860 91.385 ;
        RECT 21.530 89.775 21.870 91.215 ;
        RECT 23.655 91.065 24.695 91.215 ;
        RECT 26.520 89.775 26.860 91.215 ;
        RECT 21.530 89.605 26.860 89.775 ;
        RECT 27.290 92.950 32.620 93.120 ;
        RECT 27.290 91.385 27.630 92.950 ;
        RECT 29.415 91.385 30.455 91.525 ;
        RECT 32.280 91.385 32.620 92.950 ;
        RECT 27.290 91.215 32.620 91.385 ;
        RECT 27.290 89.775 27.630 91.215 ;
        RECT 29.415 91.065 30.455 91.215 ;
        RECT 32.280 89.775 32.620 91.215 ;
        RECT 27.290 89.605 32.620 89.775 ;
        RECT 33.050 92.950 38.380 93.120 ;
        RECT 33.050 91.385 33.390 92.950 ;
        RECT 35.175 91.385 36.215 91.525 ;
        RECT 38.040 91.385 38.380 92.950 ;
        RECT 33.050 91.215 38.380 91.385 ;
        RECT 33.050 89.775 33.390 91.215 ;
        RECT 35.175 91.065 36.215 91.215 ;
        RECT 38.040 89.775 38.380 91.215 ;
        RECT 33.050 89.605 38.380 89.775 ;
        RECT 38.810 92.950 44.140 93.120 ;
        RECT 38.810 91.385 39.150 92.950 ;
        RECT 40.935 91.385 41.975 91.525 ;
        RECT 43.800 91.385 44.140 92.950 ;
        RECT 38.810 91.215 44.140 91.385 ;
        RECT 38.810 89.775 39.150 91.215 ;
        RECT 40.935 91.065 41.975 91.215 ;
        RECT 43.800 89.775 44.140 91.215 ;
        RECT 38.810 89.605 44.140 89.775 ;
        RECT 44.570 92.950 49.900 93.120 ;
        RECT 44.570 91.385 44.910 92.950 ;
        RECT 46.695 91.385 47.735 91.525 ;
        RECT 49.560 91.385 49.900 92.950 ;
        RECT 44.570 91.215 49.900 91.385 ;
        RECT 44.570 89.775 44.910 91.215 ;
        RECT 46.695 91.065 47.735 91.215 ;
        RECT 49.560 89.775 49.900 91.215 ;
        RECT 44.570 89.605 49.900 89.775 ;
        RECT 51.905 92.890 52.075 95.130 ;
        RECT 51.905 88.350 52.745 92.890 ;
        RECT 54.155 88.350 54.325 92.890 ;
        RECT 55.735 88.350 55.905 92.890 ;
        RECT 57.315 88.350 57.485 92.890 ;
        RECT 58.895 88.350 59.065 92.890 ;
        RECT 60.475 88.350 60.645 92.890 ;
        RECT 62.055 88.350 62.225 92.890 ;
        RECT 63.635 88.350 63.805 92.890 ;
        RECT 65.215 88.350 65.385 92.890 ;
        RECT 66.795 88.350 66.965 92.890 ;
        RECT 68.375 88.350 68.545 92.890 ;
        RECT 51.905 86.125 52.075 88.350 ;
        RECT 69.835 86.125 70.005 95.130 ;
        RECT 51.905 85.955 70.005 86.125 ;
      LAYER mcon ;
        RECT 16.550 164.780 16.720 164.950 ;
        RECT 16.910 164.780 17.080 164.950 ;
        RECT 17.270 164.780 17.440 164.950 ;
        RECT 17.630 164.780 17.800 164.950 ;
        RECT 17.990 164.780 18.160 164.950 ;
        RECT 18.350 164.780 18.520 164.950 ;
        RECT 18.710 164.780 18.880 164.950 ;
        RECT 19.070 164.780 19.240 164.950 ;
        RECT 19.430 164.780 19.600 164.950 ;
        RECT 19.790 164.780 19.960 164.950 ;
        RECT 20.315 164.780 20.485 164.950 ;
        RECT 20.675 164.780 20.845 164.950 ;
        RECT 21.035 164.780 21.205 164.950 ;
        RECT 21.395 164.780 21.565 164.950 ;
        RECT 21.755 164.780 21.925 164.950 ;
        RECT 22.115 164.780 22.285 164.950 ;
        RECT 22.475 164.780 22.645 164.950 ;
        RECT 22.835 164.780 23.005 164.950 ;
        RECT 23.195 164.780 23.365 164.950 ;
        RECT 23.555 164.780 23.725 164.950 ;
        RECT 23.915 164.780 24.085 164.950 ;
        RECT 24.275 164.780 24.445 164.950 ;
        RECT 24.780 164.780 24.950 164.950 ;
        RECT 25.140 164.780 25.310 164.950 ;
        RECT 25.500 164.780 25.670 164.950 ;
        RECT 25.860 164.780 26.030 164.950 ;
        RECT 26.220 164.780 26.390 164.950 ;
        RECT 26.580 164.780 26.750 164.950 ;
        RECT 26.940 164.780 27.110 164.950 ;
        RECT 27.300 164.780 27.470 164.950 ;
        RECT 27.660 164.780 27.830 164.950 ;
        RECT 28.020 164.780 28.190 164.950 ;
        RECT 28.380 164.780 28.550 164.950 ;
        RECT 28.740 164.780 28.910 164.950 ;
        RECT 29.265 164.780 29.435 164.950 ;
        RECT 29.625 164.780 29.795 164.950 ;
        RECT 29.985 164.780 30.155 164.950 ;
        RECT 30.345 164.780 30.515 164.950 ;
        RECT 30.705 164.780 30.875 164.950 ;
        RECT 16.565 164.010 16.735 164.180 ;
        RECT 17.445 164.010 17.615 164.180 ;
        RECT 16.565 163.650 16.735 163.820 ;
        RECT 17.445 163.650 17.615 163.820 ;
        RECT 16.565 163.290 16.735 163.460 ;
        RECT 17.445 163.290 17.615 163.460 ;
        RECT 16.565 162.930 16.735 163.100 ;
        RECT 17.445 162.930 17.615 163.100 ;
        RECT 16.565 162.570 16.735 162.740 ;
        RECT 17.445 162.570 17.615 162.740 ;
        RECT 16.565 162.210 16.735 162.380 ;
        RECT 17.445 162.210 17.615 162.380 ;
        RECT 16.565 161.850 16.735 162.020 ;
        RECT 17.445 161.850 17.615 162.020 ;
        RECT 16.565 161.490 16.735 161.660 ;
        RECT 17.445 161.490 17.615 161.660 ;
        RECT 16.565 161.130 16.735 161.300 ;
        RECT 17.445 161.130 17.615 161.300 ;
        RECT 16.565 160.770 16.735 160.940 ;
        RECT 17.445 160.770 17.615 160.940 ;
        RECT 16.565 160.410 16.735 160.580 ;
        RECT 17.445 160.410 17.615 160.580 ;
        RECT 16.565 160.050 16.735 160.220 ;
        RECT 17.445 160.050 17.615 160.220 ;
        RECT 16.565 159.690 16.735 159.860 ;
        RECT 17.445 159.690 17.615 159.860 ;
        RECT 16.565 159.330 16.735 159.500 ;
        RECT 17.445 159.330 17.615 159.500 ;
        RECT 16.565 158.970 16.735 159.140 ;
        RECT 17.445 158.970 17.615 159.140 ;
        RECT 16.565 158.610 16.735 158.780 ;
        RECT 17.445 158.610 17.615 158.780 ;
        RECT 16.565 158.250 16.735 158.420 ;
        RECT 17.445 158.250 17.615 158.420 ;
        RECT 21.465 164.010 21.635 164.180 ;
        RECT 21.465 163.650 21.635 163.820 ;
        RECT 21.465 163.290 21.635 163.460 ;
        RECT 21.465 162.930 21.635 163.100 ;
        RECT 21.465 162.570 21.635 162.740 ;
        RECT 21.465 162.210 21.635 162.380 ;
        RECT 21.465 161.850 21.635 162.020 ;
        RECT 21.465 161.490 21.635 161.660 ;
        RECT 21.465 161.130 21.635 161.300 ;
        RECT 21.465 160.770 21.635 160.940 ;
        RECT 21.465 160.410 21.635 160.580 ;
        RECT 21.465 160.050 21.635 160.220 ;
        RECT 21.465 159.690 21.635 159.860 ;
        RECT 21.465 159.330 21.635 159.500 ;
        RECT 21.465 158.970 21.635 159.140 ;
        RECT 21.465 158.610 21.635 158.780 ;
        RECT 21.465 158.250 21.635 158.420 ;
        RECT 25.525 164.010 25.695 164.180 ;
        RECT 25.525 163.650 25.695 163.820 ;
        RECT 25.525 163.290 25.695 163.460 ;
        RECT 25.525 162.930 25.695 163.100 ;
        RECT 25.525 162.570 25.695 162.740 ;
        RECT 25.525 162.210 25.695 162.380 ;
        RECT 25.525 161.850 25.695 162.020 ;
        RECT 25.525 161.490 25.695 161.660 ;
        RECT 25.525 161.130 25.695 161.300 ;
        RECT 25.525 160.770 25.695 160.940 ;
        RECT 25.525 160.410 25.695 160.580 ;
        RECT 25.525 160.050 25.695 160.220 ;
        RECT 25.525 159.690 25.695 159.860 ;
        RECT 25.525 159.330 25.695 159.500 ;
        RECT 25.525 158.970 25.695 159.140 ;
        RECT 25.525 158.610 25.695 158.780 ;
        RECT 25.525 158.250 25.695 158.420 ;
        RECT 29.550 164.010 29.720 164.180 ;
        RECT 30.690 164.010 30.860 164.180 ;
        RECT 29.550 163.650 29.720 163.820 ;
        RECT 30.690 163.650 30.860 163.820 ;
        RECT 29.550 163.290 29.720 163.460 ;
        RECT 30.690 163.290 30.860 163.460 ;
        RECT 29.550 162.930 29.720 163.100 ;
        RECT 30.690 162.930 30.860 163.100 ;
        RECT 29.550 162.570 29.720 162.740 ;
        RECT 30.690 162.570 30.860 162.740 ;
        RECT 29.550 162.210 29.720 162.380 ;
        RECT 30.690 162.210 30.860 162.380 ;
        RECT 29.550 161.850 29.720 162.020 ;
        RECT 30.690 161.850 30.860 162.020 ;
        RECT 29.550 161.490 29.720 161.660 ;
        RECT 30.690 161.490 30.860 161.660 ;
        RECT 29.550 161.130 29.720 161.300 ;
        RECT 30.690 161.130 30.860 161.300 ;
        RECT 29.550 160.770 29.720 160.940 ;
        RECT 30.690 160.770 30.860 160.940 ;
        RECT 29.550 160.410 29.720 160.580 ;
        RECT 30.690 160.410 30.860 160.580 ;
        RECT 29.550 160.050 29.720 160.220 ;
        RECT 30.690 160.050 30.860 160.220 ;
        RECT 29.550 159.690 29.720 159.860 ;
        RECT 30.690 159.690 30.860 159.860 ;
        RECT 29.550 159.330 29.720 159.500 ;
        RECT 30.690 159.330 30.860 159.500 ;
        RECT 29.550 158.970 29.720 159.140 ;
        RECT 30.690 158.970 30.860 159.140 ;
        RECT 29.550 158.610 29.720 158.780 ;
        RECT 30.690 158.610 30.860 158.780 ;
        RECT 29.550 158.250 29.720 158.420 ;
        RECT 30.690 158.250 30.860 158.420 ;
        RECT 32.275 164.780 32.445 164.950 ;
        RECT 32.635 164.780 32.805 164.950 ;
        RECT 32.995 164.780 33.165 164.950 ;
        RECT 33.355 164.780 33.525 164.950 ;
        RECT 33.715 164.780 33.885 164.950 ;
        RECT 34.240 164.780 34.410 164.950 ;
        RECT 34.600 164.780 34.770 164.950 ;
        RECT 34.960 164.780 35.130 164.950 ;
        RECT 35.320 164.780 35.490 164.950 ;
        RECT 35.680 164.780 35.850 164.950 ;
        RECT 36.040 164.780 36.210 164.950 ;
        RECT 36.400 164.780 36.570 164.950 ;
        RECT 36.760 164.780 36.930 164.950 ;
        RECT 37.120 164.780 37.290 164.950 ;
        RECT 37.480 164.780 37.650 164.950 ;
        RECT 37.840 164.780 38.010 164.950 ;
        RECT 38.200 164.780 38.370 164.950 ;
        RECT 38.705 164.780 38.875 164.950 ;
        RECT 39.065 164.780 39.235 164.950 ;
        RECT 39.425 164.780 39.595 164.950 ;
        RECT 39.785 164.780 39.955 164.950 ;
        RECT 40.145 164.780 40.315 164.950 ;
        RECT 40.505 164.780 40.675 164.950 ;
        RECT 40.865 164.780 41.035 164.950 ;
        RECT 41.225 164.780 41.395 164.950 ;
        RECT 41.585 164.780 41.755 164.950 ;
        RECT 41.945 164.780 42.115 164.950 ;
        RECT 42.305 164.780 42.475 164.950 ;
        RECT 42.665 164.780 42.835 164.950 ;
        RECT 43.190 164.780 43.360 164.950 ;
        RECT 43.550 164.780 43.720 164.950 ;
        RECT 43.910 164.780 44.080 164.950 ;
        RECT 44.270 164.780 44.440 164.950 ;
        RECT 44.630 164.780 44.800 164.950 ;
        RECT 44.990 164.780 45.160 164.950 ;
        RECT 45.350 164.780 45.520 164.950 ;
        RECT 45.710 164.780 45.880 164.950 ;
        RECT 46.070 164.780 46.240 164.950 ;
        RECT 46.430 164.780 46.600 164.950 ;
        RECT 32.290 164.010 32.460 164.180 ;
        RECT 33.430 164.010 33.600 164.180 ;
        RECT 32.290 163.650 32.460 163.820 ;
        RECT 33.430 163.650 33.600 163.820 ;
        RECT 32.290 163.290 32.460 163.460 ;
        RECT 33.430 163.290 33.600 163.460 ;
        RECT 32.290 162.930 32.460 163.100 ;
        RECT 33.430 162.930 33.600 163.100 ;
        RECT 32.290 162.570 32.460 162.740 ;
        RECT 33.430 162.570 33.600 162.740 ;
        RECT 32.290 162.210 32.460 162.380 ;
        RECT 33.430 162.210 33.600 162.380 ;
        RECT 32.290 161.850 32.460 162.020 ;
        RECT 33.430 161.850 33.600 162.020 ;
        RECT 32.290 161.490 32.460 161.660 ;
        RECT 33.430 161.490 33.600 161.660 ;
        RECT 32.290 161.130 32.460 161.300 ;
        RECT 33.430 161.130 33.600 161.300 ;
        RECT 32.290 160.770 32.460 160.940 ;
        RECT 33.430 160.770 33.600 160.940 ;
        RECT 32.290 160.410 32.460 160.580 ;
        RECT 33.430 160.410 33.600 160.580 ;
        RECT 32.290 160.050 32.460 160.220 ;
        RECT 33.430 160.050 33.600 160.220 ;
        RECT 32.290 159.690 32.460 159.860 ;
        RECT 33.430 159.690 33.600 159.860 ;
        RECT 32.290 159.330 32.460 159.500 ;
        RECT 33.430 159.330 33.600 159.500 ;
        RECT 32.290 158.970 32.460 159.140 ;
        RECT 33.430 158.970 33.600 159.140 ;
        RECT 32.290 158.610 32.460 158.780 ;
        RECT 33.430 158.610 33.600 158.780 ;
        RECT 32.290 158.250 32.460 158.420 ;
        RECT 33.430 158.250 33.600 158.420 ;
        RECT 37.455 164.010 37.625 164.180 ;
        RECT 37.455 163.650 37.625 163.820 ;
        RECT 37.455 163.290 37.625 163.460 ;
        RECT 37.455 162.930 37.625 163.100 ;
        RECT 37.455 162.570 37.625 162.740 ;
        RECT 37.455 162.210 37.625 162.380 ;
        RECT 37.455 161.850 37.625 162.020 ;
        RECT 37.455 161.490 37.625 161.660 ;
        RECT 37.455 161.130 37.625 161.300 ;
        RECT 37.455 160.770 37.625 160.940 ;
        RECT 37.455 160.410 37.625 160.580 ;
        RECT 37.455 160.050 37.625 160.220 ;
        RECT 37.455 159.690 37.625 159.860 ;
        RECT 37.455 159.330 37.625 159.500 ;
        RECT 37.455 158.970 37.625 159.140 ;
        RECT 37.455 158.610 37.625 158.780 ;
        RECT 37.455 158.250 37.625 158.420 ;
        RECT 41.515 164.010 41.685 164.180 ;
        RECT 41.515 163.650 41.685 163.820 ;
        RECT 41.515 163.290 41.685 163.460 ;
        RECT 41.515 162.930 41.685 163.100 ;
        RECT 41.515 162.570 41.685 162.740 ;
        RECT 41.515 162.210 41.685 162.380 ;
        RECT 41.515 161.850 41.685 162.020 ;
        RECT 41.515 161.490 41.685 161.660 ;
        RECT 41.515 161.130 41.685 161.300 ;
        RECT 41.515 160.770 41.685 160.940 ;
        RECT 41.515 160.410 41.685 160.580 ;
        RECT 41.515 160.050 41.685 160.220 ;
        RECT 41.515 159.690 41.685 159.860 ;
        RECT 41.515 159.330 41.685 159.500 ;
        RECT 41.515 158.970 41.685 159.140 ;
        RECT 41.515 158.610 41.685 158.780 ;
        RECT 41.515 158.250 41.685 158.420 ;
        RECT 45.535 164.010 45.705 164.180 ;
        RECT 46.415 164.010 46.585 164.180 ;
        RECT 45.535 163.650 45.705 163.820 ;
        RECT 46.415 163.650 46.585 163.820 ;
        RECT 45.535 163.290 45.705 163.460 ;
        RECT 46.415 163.290 46.585 163.460 ;
        RECT 45.535 162.930 45.705 163.100 ;
        RECT 46.415 162.930 46.585 163.100 ;
        RECT 45.535 162.570 45.705 162.740 ;
        RECT 46.415 162.570 46.585 162.740 ;
        RECT 45.535 162.210 45.705 162.380 ;
        RECT 46.415 162.210 46.585 162.380 ;
        RECT 45.535 161.850 45.705 162.020 ;
        RECT 46.415 161.850 46.585 162.020 ;
        RECT 45.535 161.490 45.705 161.660 ;
        RECT 46.415 161.490 46.585 161.660 ;
        RECT 45.535 161.130 45.705 161.300 ;
        RECT 46.415 161.130 46.585 161.300 ;
        RECT 45.535 160.770 45.705 160.940 ;
        RECT 46.415 160.770 46.585 160.940 ;
        RECT 45.535 160.410 45.705 160.580 ;
        RECT 46.415 160.410 46.585 160.580 ;
        RECT 45.535 160.050 45.705 160.220 ;
        RECT 46.415 160.050 46.585 160.220 ;
        RECT 45.535 159.690 45.705 159.860 ;
        RECT 46.415 159.690 46.585 159.860 ;
        RECT 45.535 159.330 45.705 159.500 ;
        RECT 46.415 159.330 46.585 159.500 ;
        RECT 45.535 158.970 45.705 159.140 ;
        RECT 46.415 158.970 46.585 159.140 ;
        RECT 45.535 158.610 45.705 158.780 ;
        RECT 46.415 158.610 46.585 158.780 ;
        RECT 45.535 158.250 45.705 158.420 ;
        RECT 46.415 158.250 46.585 158.420 ;
        RECT 16.565 157.890 16.735 158.060 ;
        RECT 17.445 157.890 17.615 158.060 ;
        RECT 21.465 157.890 21.635 158.060 ;
        RECT 25.525 157.890 25.695 158.060 ;
        RECT 29.550 157.890 29.720 158.060 ;
        RECT 30.690 157.890 30.860 158.060 ;
        RECT 16.550 157.355 16.720 157.525 ;
        RECT 16.910 157.355 17.080 157.525 ;
        RECT 17.270 157.355 17.440 157.525 ;
        RECT 17.630 157.355 17.800 157.525 ;
        RECT 17.990 157.355 18.160 157.525 ;
        RECT 18.350 157.355 18.520 157.525 ;
        RECT 18.710 157.355 18.880 157.525 ;
        RECT 19.070 157.355 19.240 157.525 ;
        RECT 19.430 157.355 19.600 157.525 ;
        RECT 19.790 157.355 19.960 157.525 ;
        RECT 20.315 157.355 20.485 157.525 ;
        RECT 20.675 157.355 20.845 157.525 ;
        RECT 21.035 157.355 21.205 157.525 ;
        RECT 21.395 157.355 21.565 157.525 ;
        RECT 21.755 157.355 21.925 157.525 ;
        RECT 22.115 157.355 22.285 157.525 ;
        RECT 22.475 157.355 22.645 157.525 ;
        RECT 22.835 157.355 23.005 157.525 ;
        RECT 23.195 157.355 23.365 157.525 ;
        RECT 23.555 157.355 23.725 157.525 ;
        RECT 23.915 157.355 24.085 157.525 ;
        RECT 24.275 157.355 24.445 157.525 ;
        RECT 24.780 157.355 24.950 157.525 ;
        RECT 25.140 157.355 25.310 157.525 ;
        RECT 25.500 157.355 25.670 157.525 ;
        RECT 25.860 157.355 26.030 157.525 ;
        RECT 26.220 157.355 26.390 157.525 ;
        RECT 26.580 157.355 26.750 157.525 ;
        RECT 26.940 157.355 27.110 157.525 ;
        RECT 27.300 157.355 27.470 157.525 ;
        RECT 27.660 157.355 27.830 157.525 ;
        RECT 28.020 157.355 28.190 157.525 ;
        RECT 28.380 157.355 28.550 157.525 ;
        RECT 28.740 157.355 28.910 157.525 ;
        RECT 29.265 157.355 29.435 157.525 ;
        RECT 29.625 157.355 29.795 157.525 ;
        RECT 29.985 157.355 30.155 157.525 ;
        RECT 30.345 157.355 30.515 157.525 ;
        RECT 30.705 157.355 30.875 157.525 ;
        RECT 32.290 157.890 32.460 158.060 ;
        RECT 33.430 157.890 33.600 158.060 ;
        RECT 37.455 157.890 37.625 158.060 ;
        RECT 41.515 157.890 41.685 158.060 ;
        RECT 45.535 157.890 45.705 158.060 ;
        RECT 46.415 157.890 46.585 158.060 ;
        RECT 32.275 157.355 32.445 157.525 ;
        RECT 32.635 157.355 32.805 157.525 ;
        RECT 32.995 157.355 33.165 157.525 ;
        RECT 33.355 157.355 33.525 157.525 ;
        RECT 33.715 157.355 33.885 157.525 ;
        RECT 34.240 157.355 34.410 157.525 ;
        RECT 34.600 157.355 34.770 157.525 ;
        RECT 34.960 157.355 35.130 157.525 ;
        RECT 35.320 157.355 35.490 157.525 ;
        RECT 35.680 157.355 35.850 157.525 ;
        RECT 36.040 157.355 36.210 157.525 ;
        RECT 36.400 157.355 36.570 157.525 ;
        RECT 36.760 157.355 36.930 157.525 ;
        RECT 37.120 157.355 37.290 157.525 ;
        RECT 37.480 157.355 37.650 157.525 ;
        RECT 37.840 157.355 38.010 157.525 ;
        RECT 38.200 157.355 38.370 157.525 ;
        RECT 38.705 157.355 38.875 157.525 ;
        RECT 39.065 157.355 39.235 157.525 ;
        RECT 39.425 157.355 39.595 157.525 ;
        RECT 39.785 157.355 39.955 157.525 ;
        RECT 40.145 157.355 40.315 157.525 ;
        RECT 40.505 157.355 40.675 157.525 ;
        RECT 40.865 157.355 41.035 157.525 ;
        RECT 41.225 157.355 41.395 157.525 ;
        RECT 41.585 157.355 41.755 157.525 ;
        RECT 41.945 157.355 42.115 157.525 ;
        RECT 42.305 157.355 42.475 157.525 ;
        RECT 42.665 157.355 42.835 157.525 ;
        RECT 43.190 157.355 43.360 157.525 ;
        RECT 43.550 157.355 43.720 157.525 ;
        RECT 43.910 157.355 44.080 157.525 ;
        RECT 44.270 157.355 44.440 157.525 ;
        RECT 44.630 157.355 44.800 157.525 ;
        RECT 44.990 157.355 45.160 157.525 ;
        RECT 45.350 157.355 45.520 157.525 ;
        RECT 45.710 157.355 45.880 157.525 ;
        RECT 46.070 157.355 46.240 157.525 ;
        RECT 46.430 157.355 46.600 157.525 ;
        RECT 53.980 113.740 54.150 113.910 ;
        RECT 54.650 113.740 54.820 113.910 ;
        RECT 53.980 113.380 54.150 113.550 ;
        RECT 54.650 113.380 54.820 113.550 ;
        RECT 53.980 113.020 54.150 113.190 ;
        RECT 54.650 113.020 54.820 113.190 ;
        RECT 53.980 112.660 54.150 112.830 ;
        RECT 54.650 112.660 54.820 112.830 ;
        RECT 56.230 113.740 56.400 113.910 ;
        RECT 56.230 113.380 56.400 113.550 ;
        RECT 56.230 113.020 56.400 113.190 ;
        RECT 56.230 112.660 56.400 112.830 ;
        RECT 57.810 113.740 57.980 113.910 ;
        RECT 57.810 113.380 57.980 113.550 ;
        RECT 57.810 113.020 57.980 113.190 ;
        RECT 57.810 112.660 57.980 112.830 ;
        RECT 59.390 113.740 59.560 113.910 ;
        RECT 60.060 113.740 60.230 113.910 ;
        RECT 59.390 113.380 59.560 113.550 ;
        RECT 60.060 113.380 60.230 113.550 ;
        RECT 59.390 113.020 59.560 113.190 ;
        RECT 60.060 113.020 60.230 113.190 ;
        RECT 59.390 112.660 59.560 112.830 ;
        RECT 60.060 112.660 60.230 112.830 ;
        RECT 61.910 113.740 62.080 113.910 ;
        RECT 62.580 113.740 62.750 113.910 ;
        RECT 61.910 113.380 62.080 113.550 ;
        RECT 62.580 113.380 62.750 113.550 ;
        RECT 61.910 113.020 62.080 113.190 ;
        RECT 62.580 113.020 62.750 113.190 ;
        RECT 61.910 112.660 62.080 112.830 ;
        RECT 62.580 112.660 62.750 112.830 ;
        RECT 64.160 113.740 64.330 113.910 ;
        RECT 64.160 113.380 64.330 113.550 ;
        RECT 64.160 113.020 64.330 113.190 ;
        RECT 64.160 112.660 64.330 112.830 ;
        RECT 65.740 113.740 65.910 113.910 ;
        RECT 65.740 113.380 65.910 113.550 ;
        RECT 65.740 113.020 65.910 113.190 ;
        RECT 65.740 112.660 65.910 112.830 ;
        RECT 67.320 113.740 67.490 113.910 ;
        RECT 67.320 113.380 67.490 113.550 ;
        RECT 67.320 113.020 67.490 113.190 ;
        RECT 67.320 112.660 67.490 112.830 ;
        RECT 68.900 113.740 69.070 113.910 ;
        RECT 68.900 113.380 69.070 113.550 ;
        RECT 68.900 113.020 69.070 113.190 ;
        RECT 68.900 112.660 69.070 112.830 ;
        RECT 70.360 113.740 70.530 113.910 ;
        RECT 70.360 113.380 70.530 113.550 ;
        RECT 70.360 113.020 70.530 113.190 ;
        RECT 70.360 112.660 70.530 112.830 ;
        RECT 15.455 102.390 15.625 102.560 ;
        RECT 15.815 102.390 15.985 102.560 ;
        RECT 16.835 102.390 17.005 102.560 ;
        RECT 17.195 102.390 17.365 102.560 ;
        RECT 17.555 102.390 17.725 102.560 ;
        RECT 18.745 102.390 18.915 102.560 ;
        RECT 19.270 102.420 19.440 102.590 ;
        RECT 19.630 102.420 19.800 102.590 ;
        RECT 20.575 102.420 20.745 102.590 ;
        RECT 20.935 102.420 21.105 102.590 ;
        RECT 21.295 102.420 21.465 102.590 ;
        RECT 22.135 102.420 22.305 102.590 ;
        RECT 22.495 102.420 22.665 102.590 ;
        RECT 22.855 102.420 23.025 102.590 ;
        RECT 23.695 102.420 23.865 102.590 ;
        RECT 24.055 102.420 24.225 102.590 ;
        RECT 24.415 102.420 24.585 102.590 ;
        RECT 25.255 102.420 25.425 102.590 ;
        RECT 25.615 102.420 25.785 102.590 ;
        RECT 25.975 102.420 26.145 102.590 ;
        RECT 26.815 102.420 26.985 102.590 ;
        RECT 27.175 102.420 27.345 102.590 ;
        RECT 27.535 102.420 27.705 102.590 ;
        RECT 28.375 102.420 28.545 102.590 ;
        RECT 28.735 102.420 28.905 102.590 ;
        RECT 29.095 102.420 29.265 102.590 ;
        RECT 29.935 102.420 30.105 102.590 ;
        RECT 30.295 102.420 30.465 102.590 ;
        RECT 30.655 102.420 30.825 102.590 ;
        RECT 31.540 102.420 31.710 102.590 ;
        RECT 31.900 102.420 32.070 102.590 ;
        RECT 32.735 102.390 32.905 102.560 ;
        RECT 33.095 102.390 33.265 102.560 ;
        RECT 34.115 102.390 34.285 102.560 ;
        RECT 34.475 102.390 34.645 102.560 ;
        RECT 34.835 102.390 35.005 102.560 ;
        RECT 36.025 102.390 36.195 102.560 ;
        RECT 36.550 102.420 36.720 102.590 ;
        RECT 36.910 102.420 37.080 102.590 ;
        RECT 37.855 102.420 38.025 102.590 ;
        RECT 38.215 102.420 38.385 102.590 ;
        RECT 38.575 102.420 38.745 102.590 ;
        RECT 39.415 102.420 39.585 102.590 ;
        RECT 39.775 102.420 39.945 102.590 ;
        RECT 40.135 102.420 40.305 102.590 ;
        RECT 40.975 102.420 41.145 102.590 ;
        RECT 41.335 102.420 41.505 102.590 ;
        RECT 41.695 102.420 41.865 102.590 ;
        RECT 42.535 102.420 42.705 102.590 ;
        RECT 42.895 102.420 43.065 102.590 ;
        RECT 43.255 102.420 43.425 102.590 ;
        RECT 44.095 102.420 44.265 102.590 ;
        RECT 44.455 102.420 44.625 102.590 ;
        RECT 44.815 102.420 44.985 102.590 ;
        RECT 45.655 102.420 45.825 102.590 ;
        RECT 46.015 102.420 46.185 102.590 ;
        RECT 46.375 102.420 46.545 102.590 ;
        RECT 47.215 102.420 47.385 102.590 ;
        RECT 47.575 102.420 47.745 102.590 ;
        RECT 47.935 102.420 48.105 102.590 ;
        RECT 48.820 102.420 48.990 102.590 ;
        RECT 49.180 102.420 49.350 102.590 ;
        RECT 50.015 102.390 50.185 102.560 ;
        RECT 50.375 102.390 50.545 102.560 ;
        RECT 51.395 102.390 51.565 102.560 ;
        RECT 51.755 102.390 51.925 102.560 ;
        RECT 52.115 102.390 52.285 102.560 ;
        RECT 53.305 102.390 53.475 102.560 ;
        RECT 53.830 102.420 54.000 102.590 ;
        RECT 54.190 102.420 54.360 102.590 ;
        RECT 55.135 102.420 55.305 102.590 ;
        RECT 55.495 102.420 55.665 102.590 ;
        RECT 55.855 102.420 56.025 102.590 ;
        RECT 56.695 102.420 56.865 102.590 ;
        RECT 57.055 102.420 57.225 102.590 ;
        RECT 57.415 102.420 57.585 102.590 ;
        RECT 58.255 102.420 58.425 102.590 ;
        RECT 58.615 102.420 58.785 102.590 ;
        RECT 58.975 102.420 59.145 102.590 ;
        RECT 59.815 102.420 59.985 102.590 ;
        RECT 60.175 102.420 60.345 102.590 ;
        RECT 60.535 102.420 60.705 102.590 ;
        RECT 61.375 102.420 61.545 102.590 ;
        RECT 61.735 102.420 61.905 102.590 ;
        RECT 62.095 102.420 62.265 102.590 ;
        RECT 62.935 102.420 63.105 102.590 ;
        RECT 63.295 102.420 63.465 102.590 ;
        RECT 63.655 102.420 63.825 102.590 ;
        RECT 64.495 102.420 64.665 102.590 ;
        RECT 64.855 102.420 65.025 102.590 ;
        RECT 65.215 102.420 65.385 102.590 ;
        RECT 66.100 102.420 66.270 102.590 ;
        RECT 66.460 102.420 66.630 102.590 ;
        RECT 15.490 101.910 15.660 102.080 ;
        RECT 15.970 101.910 16.140 102.080 ;
        RECT 16.450 101.910 16.620 102.080 ;
        RECT 16.930 101.910 17.100 102.080 ;
        RECT 17.410 101.910 17.580 102.080 ;
        RECT 17.890 101.910 18.060 102.080 ;
        RECT 18.370 101.910 18.540 102.080 ;
        RECT 18.850 101.910 19.020 102.080 ;
        RECT 19.330 101.910 19.500 102.080 ;
        RECT 19.810 101.910 19.980 102.080 ;
        RECT 20.290 101.910 20.460 102.080 ;
        RECT 20.770 101.910 20.940 102.080 ;
        RECT 21.250 101.910 21.420 102.080 ;
        RECT 21.730 101.910 21.900 102.080 ;
        RECT 22.210 101.910 22.380 102.080 ;
        RECT 22.690 101.910 22.860 102.080 ;
        RECT 23.170 101.910 23.340 102.080 ;
        RECT 23.650 101.910 23.820 102.080 ;
        RECT 24.130 101.910 24.300 102.080 ;
        RECT 24.610 101.910 24.780 102.080 ;
        RECT 25.090 101.910 25.260 102.080 ;
        RECT 25.570 101.910 25.740 102.080 ;
        RECT 26.050 101.910 26.220 102.080 ;
        RECT 26.530 101.910 26.700 102.080 ;
        RECT 27.010 101.910 27.180 102.080 ;
        RECT 27.490 101.910 27.660 102.080 ;
        RECT 27.970 101.910 28.140 102.080 ;
        RECT 28.450 101.910 28.620 102.080 ;
        RECT 28.930 101.910 29.100 102.080 ;
        RECT 29.410 101.910 29.580 102.080 ;
        RECT 29.890 101.910 30.060 102.080 ;
        RECT 30.370 101.910 30.540 102.080 ;
        RECT 30.850 101.910 31.020 102.080 ;
        RECT 31.330 101.910 31.500 102.080 ;
        RECT 31.810 101.910 31.980 102.080 ;
        RECT 32.290 101.910 32.460 102.080 ;
        RECT 32.770 101.910 32.940 102.080 ;
        RECT 33.250 101.910 33.420 102.080 ;
        RECT 33.730 101.910 33.900 102.080 ;
        RECT 34.210 101.910 34.380 102.080 ;
        RECT 34.690 101.910 34.860 102.080 ;
        RECT 35.170 101.910 35.340 102.080 ;
        RECT 35.650 101.910 35.820 102.080 ;
        RECT 36.130 101.910 36.300 102.080 ;
        RECT 36.610 101.910 36.780 102.080 ;
        RECT 37.090 101.910 37.260 102.080 ;
        RECT 37.570 101.910 37.740 102.080 ;
        RECT 38.050 101.910 38.220 102.080 ;
        RECT 38.530 101.910 38.700 102.080 ;
        RECT 39.010 101.910 39.180 102.080 ;
        RECT 39.490 101.910 39.660 102.080 ;
        RECT 39.970 101.910 40.140 102.080 ;
        RECT 40.450 101.910 40.620 102.080 ;
        RECT 40.930 101.910 41.100 102.080 ;
        RECT 41.410 101.910 41.580 102.080 ;
        RECT 41.890 101.910 42.060 102.080 ;
        RECT 42.370 101.910 42.540 102.080 ;
        RECT 42.850 101.910 43.020 102.080 ;
        RECT 43.330 101.910 43.500 102.080 ;
        RECT 43.810 101.910 43.980 102.080 ;
        RECT 44.290 101.910 44.460 102.080 ;
        RECT 44.770 101.910 44.940 102.080 ;
        RECT 45.250 101.910 45.420 102.080 ;
        RECT 45.730 101.910 45.900 102.080 ;
        RECT 46.210 101.910 46.380 102.080 ;
        RECT 46.690 101.910 46.860 102.080 ;
        RECT 47.170 101.910 47.340 102.080 ;
        RECT 47.650 101.910 47.820 102.080 ;
        RECT 48.130 101.910 48.300 102.080 ;
        RECT 48.610 101.910 48.780 102.080 ;
        RECT 49.090 101.910 49.260 102.080 ;
        RECT 49.570 101.910 49.740 102.080 ;
        RECT 50.050 101.910 50.220 102.080 ;
        RECT 50.530 101.910 50.700 102.080 ;
        RECT 51.010 101.910 51.180 102.080 ;
        RECT 51.490 101.910 51.660 102.080 ;
        RECT 51.970 101.910 52.140 102.080 ;
        RECT 52.450 101.910 52.620 102.080 ;
        RECT 52.930 101.910 53.100 102.080 ;
        RECT 53.410 101.910 53.580 102.080 ;
        RECT 53.890 101.910 54.060 102.080 ;
        RECT 54.370 101.910 54.540 102.080 ;
        RECT 54.850 101.910 55.020 102.080 ;
        RECT 55.330 101.910 55.500 102.080 ;
        RECT 55.810 101.910 55.980 102.080 ;
        RECT 56.290 101.910 56.460 102.080 ;
        RECT 56.770 101.910 56.940 102.080 ;
        RECT 57.250 101.910 57.420 102.080 ;
        RECT 57.730 101.910 57.900 102.080 ;
        RECT 58.210 101.910 58.380 102.080 ;
        RECT 58.690 101.910 58.860 102.080 ;
        RECT 59.170 101.910 59.340 102.080 ;
        RECT 59.650 101.910 59.820 102.080 ;
        RECT 60.130 101.910 60.300 102.080 ;
        RECT 60.610 101.910 60.780 102.080 ;
        RECT 61.090 101.910 61.260 102.080 ;
        RECT 61.570 101.910 61.740 102.080 ;
        RECT 62.050 101.910 62.220 102.080 ;
        RECT 62.530 101.910 62.700 102.080 ;
        RECT 63.010 101.910 63.180 102.080 ;
        RECT 63.490 101.910 63.660 102.080 ;
        RECT 63.970 101.910 64.140 102.080 ;
        RECT 64.450 101.910 64.620 102.080 ;
        RECT 64.930 101.910 65.100 102.080 ;
        RECT 65.410 101.910 65.580 102.080 ;
        RECT 65.890 101.910 66.060 102.080 ;
        RECT 66.370 101.910 66.540 102.080 ;
        RECT 66.850 101.910 67.020 102.080 ;
        RECT 15.455 101.430 15.625 101.600 ;
        RECT 15.815 101.430 15.985 101.600 ;
        RECT 16.835 101.430 17.005 101.600 ;
        RECT 17.195 101.430 17.365 101.600 ;
        RECT 17.555 101.430 17.725 101.600 ;
        RECT 18.745 101.430 18.915 101.600 ;
        RECT 19.270 101.400 19.440 101.570 ;
        RECT 19.630 101.400 19.800 101.570 ;
        RECT 20.575 101.400 20.745 101.570 ;
        RECT 20.935 101.400 21.105 101.570 ;
        RECT 21.295 101.400 21.465 101.570 ;
        RECT 22.135 101.400 22.305 101.570 ;
        RECT 22.495 101.400 22.665 101.570 ;
        RECT 22.855 101.400 23.025 101.570 ;
        RECT 23.695 101.400 23.865 101.570 ;
        RECT 24.055 101.400 24.225 101.570 ;
        RECT 24.415 101.400 24.585 101.570 ;
        RECT 25.255 101.400 25.425 101.570 ;
        RECT 25.615 101.400 25.785 101.570 ;
        RECT 25.975 101.400 26.145 101.570 ;
        RECT 26.815 101.400 26.985 101.570 ;
        RECT 27.175 101.400 27.345 101.570 ;
        RECT 27.535 101.400 27.705 101.570 ;
        RECT 28.375 101.400 28.545 101.570 ;
        RECT 28.735 101.400 28.905 101.570 ;
        RECT 29.095 101.400 29.265 101.570 ;
        RECT 29.935 101.400 30.105 101.570 ;
        RECT 30.295 101.400 30.465 101.570 ;
        RECT 30.655 101.400 30.825 101.570 ;
        RECT 31.540 101.400 31.710 101.570 ;
        RECT 31.900 101.400 32.070 101.570 ;
        RECT 32.735 101.430 32.905 101.600 ;
        RECT 33.095 101.430 33.265 101.600 ;
        RECT 34.115 101.430 34.285 101.600 ;
        RECT 34.475 101.430 34.645 101.600 ;
        RECT 34.835 101.430 35.005 101.600 ;
        RECT 36.025 101.430 36.195 101.600 ;
        RECT 36.550 101.400 36.720 101.570 ;
        RECT 36.910 101.400 37.080 101.570 ;
        RECT 37.855 101.400 38.025 101.570 ;
        RECT 38.215 101.400 38.385 101.570 ;
        RECT 38.575 101.400 38.745 101.570 ;
        RECT 39.415 101.400 39.585 101.570 ;
        RECT 39.775 101.400 39.945 101.570 ;
        RECT 40.135 101.400 40.305 101.570 ;
        RECT 40.975 101.400 41.145 101.570 ;
        RECT 41.335 101.400 41.505 101.570 ;
        RECT 41.695 101.400 41.865 101.570 ;
        RECT 42.535 101.400 42.705 101.570 ;
        RECT 42.895 101.400 43.065 101.570 ;
        RECT 43.255 101.400 43.425 101.570 ;
        RECT 44.095 101.400 44.265 101.570 ;
        RECT 44.455 101.400 44.625 101.570 ;
        RECT 44.815 101.400 44.985 101.570 ;
        RECT 45.655 101.400 45.825 101.570 ;
        RECT 46.015 101.400 46.185 101.570 ;
        RECT 46.375 101.400 46.545 101.570 ;
        RECT 47.215 101.400 47.385 101.570 ;
        RECT 47.575 101.400 47.745 101.570 ;
        RECT 47.935 101.400 48.105 101.570 ;
        RECT 48.820 101.400 48.990 101.570 ;
        RECT 49.180 101.400 49.350 101.570 ;
        RECT 50.015 101.430 50.185 101.600 ;
        RECT 50.375 101.430 50.545 101.600 ;
        RECT 51.395 101.430 51.565 101.600 ;
        RECT 51.755 101.430 51.925 101.600 ;
        RECT 52.115 101.430 52.285 101.600 ;
        RECT 53.305 101.430 53.475 101.600 ;
        RECT 53.830 101.400 54.000 101.570 ;
        RECT 54.190 101.400 54.360 101.570 ;
        RECT 55.135 101.400 55.305 101.570 ;
        RECT 55.495 101.400 55.665 101.570 ;
        RECT 55.855 101.400 56.025 101.570 ;
        RECT 56.695 101.400 56.865 101.570 ;
        RECT 57.055 101.400 57.225 101.570 ;
        RECT 57.415 101.400 57.585 101.570 ;
        RECT 58.255 101.400 58.425 101.570 ;
        RECT 58.615 101.400 58.785 101.570 ;
        RECT 58.975 101.400 59.145 101.570 ;
        RECT 59.815 101.400 59.985 101.570 ;
        RECT 60.175 101.400 60.345 101.570 ;
        RECT 60.535 101.400 60.705 101.570 ;
        RECT 61.375 101.400 61.545 101.570 ;
        RECT 61.735 101.400 61.905 101.570 ;
        RECT 62.095 101.400 62.265 101.570 ;
        RECT 62.935 101.400 63.105 101.570 ;
        RECT 63.295 101.400 63.465 101.570 ;
        RECT 63.655 101.400 63.825 101.570 ;
        RECT 64.495 101.400 64.665 101.570 ;
        RECT 64.855 101.400 65.025 101.570 ;
        RECT 65.215 101.400 65.385 101.570 ;
        RECT 66.100 101.400 66.270 101.570 ;
        RECT 66.460 101.400 66.630 101.570 ;
        RECT 15.870 91.210 16.040 91.380 ;
        RECT 18.270 91.210 18.440 91.380 ;
        RECT 18.630 91.210 18.800 91.380 ;
        RECT 20.835 91.210 21.005 91.380 ;
        RECT 21.630 91.210 21.800 91.380 ;
        RECT 24.030 91.210 24.200 91.380 ;
        RECT 24.390 91.210 24.560 91.380 ;
        RECT 26.595 91.210 26.765 91.380 ;
        RECT 27.390 91.210 27.560 91.380 ;
        RECT 29.790 91.210 29.960 91.380 ;
        RECT 30.150 91.210 30.320 91.380 ;
        RECT 32.355 91.210 32.525 91.380 ;
        RECT 33.150 91.210 33.320 91.380 ;
        RECT 35.550 91.210 35.720 91.380 ;
        RECT 35.910 91.210 36.080 91.380 ;
        RECT 38.115 91.210 38.285 91.380 ;
        RECT 38.910 91.210 39.080 91.380 ;
        RECT 41.310 91.210 41.480 91.380 ;
        RECT 41.670 91.210 41.840 91.380 ;
        RECT 43.875 91.210 44.045 91.380 ;
        RECT 44.670 91.210 44.840 91.380 ;
        RECT 47.070 91.210 47.240 91.380 ;
        RECT 47.430 91.210 47.600 91.380 ;
        RECT 49.635 91.210 49.805 91.380 ;
        RECT 51.905 92.515 52.075 92.685 ;
        RECT 52.575 92.515 52.745 92.685 ;
        RECT 51.905 92.155 52.075 92.325 ;
        RECT 52.575 92.155 52.745 92.325 ;
        RECT 51.905 91.795 52.075 91.965 ;
        RECT 52.575 91.795 52.745 91.965 ;
        RECT 51.905 91.435 52.075 91.605 ;
        RECT 52.575 91.435 52.745 91.605 ;
        RECT 54.155 92.515 54.325 92.685 ;
        RECT 54.155 92.155 54.325 92.325 ;
        RECT 54.155 91.795 54.325 91.965 ;
        RECT 54.155 91.435 54.325 91.605 ;
        RECT 55.735 92.515 55.905 92.685 ;
        RECT 55.735 92.155 55.905 92.325 ;
        RECT 55.735 91.795 55.905 91.965 ;
        RECT 55.735 91.435 55.905 91.605 ;
        RECT 57.315 92.515 57.485 92.685 ;
        RECT 57.315 92.155 57.485 92.325 ;
        RECT 57.315 91.795 57.485 91.965 ;
        RECT 57.315 91.435 57.485 91.605 ;
        RECT 58.895 92.515 59.065 92.685 ;
        RECT 58.895 92.155 59.065 92.325 ;
        RECT 58.895 91.795 59.065 91.965 ;
        RECT 58.895 91.435 59.065 91.605 ;
        RECT 60.475 92.515 60.645 92.685 ;
        RECT 60.475 92.155 60.645 92.325 ;
        RECT 60.475 91.795 60.645 91.965 ;
        RECT 60.475 91.435 60.645 91.605 ;
        RECT 62.055 92.515 62.225 92.685 ;
        RECT 62.055 92.155 62.225 92.325 ;
        RECT 62.055 91.795 62.225 91.965 ;
        RECT 62.055 91.435 62.225 91.605 ;
        RECT 63.635 92.515 63.805 92.685 ;
        RECT 63.635 92.155 63.805 92.325 ;
        RECT 63.635 91.795 63.805 91.965 ;
        RECT 63.635 91.435 63.805 91.605 ;
        RECT 65.215 92.515 65.385 92.685 ;
        RECT 65.215 92.155 65.385 92.325 ;
        RECT 65.215 91.795 65.385 91.965 ;
        RECT 65.215 91.435 65.385 91.605 ;
        RECT 66.795 92.515 66.965 92.685 ;
        RECT 66.795 92.155 66.965 92.325 ;
        RECT 66.795 91.795 66.965 91.965 ;
        RECT 66.795 91.435 66.965 91.605 ;
        RECT 68.375 92.515 68.545 92.685 ;
        RECT 68.375 92.155 68.545 92.325 ;
        RECT 68.375 91.795 68.545 91.965 ;
        RECT 68.375 91.435 68.545 91.605 ;
        RECT 69.835 92.515 70.005 92.685 ;
        RECT 69.835 92.155 70.005 92.325 ;
        RECT 69.835 91.795 70.005 91.965 ;
        RECT 69.835 91.435 70.005 91.605 ;
      LAYER met1 ;
        RECT 16.090 164.250 47.060 165.495 ;
        RECT 16.090 158.225 18.015 164.250 ;
        RECT 20.990 158.225 22.125 164.250 ;
        RECT 25.040 158.225 26.175 164.250 ;
        RECT 29.210 158.225 31.135 164.250 ;
        RECT 32.015 158.225 33.940 164.250 ;
        RECT 36.975 158.225 38.110 164.250 ;
        RECT 41.025 158.225 42.160 164.250 ;
        RECT 45.135 158.225 47.060 164.250 ;
        RECT 16.090 156.980 47.060 158.225 ;
        RECT 53.815 112.475 70.735 114.180 ;
        RECT 5.300 101.370 67.680 102.620 ;
        RECT 6.015 91.115 50.420 91.470 ;
        RECT 51.740 91.165 70.210 92.870 ;
        RECT 0.000 47.205 88.240 81.515 ;
      LAYER via ;
        RECT 16.565 164.825 16.825 165.085 ;
        RECT 16.905 164.825 17.165 165.085 ;
        RECT 17.225 164.825 17.485 165.085 ;
        RECT 16.565 164.500 16.825 164.760 ;
        RECT 16.905 164.500 17.165 164.760 ;
        RECT 17.225 164.500 17.485 164.760 ;
        RECT 16.565 164.170 16.825 164.430 ;
        RECT 16.905 164.170 17.165 164.430 ;
        RECT 17.225 164.170 17.485 164.430 ;
        RECT 16.565 163.680 16.825 163.940 ;
        RECT 16.905 163.680 17.165 163.940 ;
        RECT 17.225 163.680 17.485 163.940 ;
        RECT 16.565 163.355 16.825 163.615 ;
        RECT 16.905 163.355 17.165 163.615 ;
        RECT 17.225 163.355 17.485 163.615 ;
        RECT 16.565 163.025 16.825 163.285 ;
        RECT 16.905 163.025 17.165 163.285 ;
        RECT 17.225 163.025 17.485 163.285 ;
        RECT 16.565 162.620 16.825 162.880 ;
        RECT 16.905 162.620 17.165 162.880 ;
        RECT 17.225 162.620 17.485 162.880 ;
        RECT 16.565 162.295 16.825 162.555 ;
        RECT 16.905 162.295 17.165 162.555 ;
        RECT 17.225 162.295 17.485 162.555 ;
        RECT 16.565 161.965 16.825 162.225 ;
        RECT 16.905 161.965 17.165 162.225 ;
        RECT 17.225 161.965 17.485 162.225 ;
        RECT 16.565 161.475 16.825 161.735 ;
        RECT 16.905 161.475 17.165 161.735 ;
        RECT 17.225 161.475 17.485 161.735 ;
        RECT 16.565 161.150 16.825 161.410 ;
        RECT 16.905 161.150 17.165 161.410 ;
        RECT 17.225 161.150 17.485 161.410 ;
        RECT 16.565 160.820 16.825 161.080 ;
        RECT 16.905 160.820 17.165 161.080 ;
        RECT 17.225 160.820 17.485 161.080 ;
        RECT 16.565 160.315 16.825 160.575 ;
        RECT 16.905 160.315 17.165 160.575 ;
        RECT 17.225 160.315 17.485 160.575 ;
        RECT 16.565 159.990 16.825 160.250 ;
        RECT 16.905 159.990 17.165 160.250 ;
        RECT 17.225 159.990 17.485 160.250 ;
        RECT 16.565 159.660 16.825 159.920 ;
        RECT 16.905 159.660 17.165 159.920 ;
        RECT 17.225 159.660 17.485 159.920 ;
        RECT 16.565 159.170 16.825 159.430 ;
        RECT 16.905 159.170 17.165 159.430 ;
        RECT 17.225 159.170 17.485 159.430 ;
        RECT 16.565 158.845 16.825 159.105 ;
        RECT 16.905 158.845 17.165 159.105 ;
        RECT 17.225 158.845 17.485 159.105 ;
        RECT 16.565 158.515 16.825 158.775 ;
        RECT 16.905 158.515 17.165 158.775 ;
        RECT 17.225 158.515 17.485 158.775 ;
        RECT 16.565 158.110 16.825 158.370 ;
        RECT 16.905 158.110 17.165 158.370 ;
        RECT 17.225 158.110 17.485 158.370 ;
        RECT 16.565 157.785 16.825 158.045 ;
        RECT 16.905 157.785 17.165 158.045 ;
        RECT 17.225 157.785 17.485 158.045 ;
        RECT 16.565 157.455 16.825 157.715 ;
        RECT 16.905 157.455 17.165 157.715 ;
        RECT 17.225 157.455 17.485 157.715 ;
        RECT 63.215 113.755 63.475 114.015 ;
        RECT 63.555 113.755 63.815 114.015 ;
        RECT 64.120 113.755 64.380 114.015 ;
        RECT 64.460 113.755 64.720 114.015 ;
        RECT 64.780 113.755 65.040 114.015 ;
        RECT 65.185 113.755 65.445 114.015 ;
        RECT 65.525 113.755 65.785 114.015 ;
        RECT 65.845 113.755 66.105 114.015 ;
        RECT 66.330 113.755 66.590 114.015 ;
        RECT 63.215 113.430 63.475 113.690 ;
        RECT 63.555 113.430 63.815 113.690 ;
        RECT 64.120 113.430 64.380 113.690 ;
        RECT 64.460 113.430 64.720 113.690 ;
        RECT 64.780 113.430 65.040 113.690 ;
        RECT 65.185 113.430 65.445 113.690 ;
        RECT 65.525 113.430 65.785 113.690 ;
        RECT 65.845 113.430 66.105 113.690 ;
        RECT 66.330 113.430 66.590 113.690 ;
        RECT 63.215 113.005 63.475 113.265 ;
        RECT 63.555 113.005 63.815 113.265 ;
        RECT 64.120 113.005 64.380 113.265 ;
        RECT 64.460 113.005 64.720 113.265 ;
        RECT 64.780 113.005 65.040 113.265 ;
        RECT 65.185 113.005 65.445 113.265 ;
        RECT 65.525 113.005 65.785 113.265 ;
        RECT 65.845 113.005 66.105 113.265 ;
        RECT 66.330 113.005 66.590 113.265 ;
        RECT 63.215 112.680 63.475 112.940 ;
        RECT 63.555 112.680 63.815 112.940 ;
        RECT 64.120 112.680 64.380 112.940 ;
        RECT 64.460 112.680 64.720 112.940 ;
        RECT 64.780 112.680 65.040 112.940 ;
        RECT 65.185 112.680 65.445 112.940 ;
        RECT 65.525 112.680 65.785 112.940 ;
        RECT 65.845 112.680 66.105 112.940 ;
        RECT 66.330 112.680 66.590 112.940 ;
        RECT 6.145 102.160 6.405 102.420 ;
        RECT 6.485 102.160 6.745 102.420 ;
        RECT 6.805 102.160 7.065 102.420 ;
        RECT 7.210 102.160 7.470 102.420 ;
        RECT 7.550 102.160 7.810 102.420 ;
        RECT 8.000 102.160 8.260 102.420 ;
        RECT 8.340 102.160 8.600 102.420 ;
        RECT 8.660 102.160 8.920 102.420 ;
        RECT 9.065 102.160 9.325 102.420 ;
        RECT 9.405 102.160 9.665 102.420 ;
        RECT 6.145 101.835 6.405 102.095 ;
        RECT 6.485 101.835 6.745 102.095 ;
        RECT 6.805 101.835 7.065 102.095 ;
        RECT 7.210 101.835 7.470 102.095 ;
        RECT 7.550 101.835 7.810 102.095 ;
        RECT 8.000 101.835 8.260 102.095 ;
        RECT 8.340 101.835 8.600 102.095 ;
        RECT 8.660 101.835 8.920 102.095 ;
        RECT 9.065 101.835 9.325 102.095 ;
        RECT 9.405 101.835 9.665 102.095 ;
        RECT 6.145 101.505 6.405 101.765 ;
        RECT 6.485 101.505 6.745 101.765 ;
        RECT 6.805 101.505 7.065 101.765 ;
        RECT 7.210 101.505 7.470 101.765 ;
        RECT 7.550 101.505 7.810 101.765 ;
        RECT 8.000 101.505 8.260 101.765 ;
        RECT 8.340 101.505 8.600 101.765 ;
        RECT 8.660 101.505 8.920 101.765 ;
        RECT 9.065 101.505 9.325 101.765 ;
        RECT 9.405 101.505 9.665 101.765 ;
        RECT 62.945 92.435 63.205 92.695 ;
        RECT 63.285 92.435 63.545 92.695 ;
        RECT 63.850 92.435 64.110 92.695 ;
        RECT 64.190 92.435 64.450 92.695 ;
        RECT 64.510 92.435 64.770 92.695 ;
        RECT 64.915 92.435 65.175 92.695 ;
        RECT 65.255 92.435 65.515 92.695 ;
        RECT 65.575 92.435 65.835 92.695 ;
        RECT 66.060 92.435 66.320 92.695 ;
        RECT 62.945 92.110 63.205 92.370 ;
        RECT 63.285 92.110 63.545 92.370 ;
        RECT 63.850 92.110 64.110 92.370 ;
        RECT 64.190 92.110 64.450 92.370 ;
        RECT 64.510 92.110 64.770 92.370 ;
        RECT 64.915 92.110 65.175 92.370 ;
        RECT 65.255 92.110 65.515 92.370 ;
        RECT 65.575 92.110 65.835 92.370 ;
        RECT 66.060 92.110 66.320 92.370 ;
        RECT 62.945 91.685 63.205 91.945 ;
        RECT 63.285 91.685 63.545 91.945 ;
        RECT 63.850 91.685 64.110 91.945 ;
        RECT 64.190 91.685 64.450 91.945 ;
        RECT 64.510 91.685 64.770 91.945 ;
        RECT 64.915 91.685 65.175 91.945 ;
        RECT 65.255 91.685 65.515 91.945 ;
        RECT 65.575 91.685 65.835 91.945 ;
        RECT 66.060 91.685 66.320 91.945 ;
        RECT 6.395 91.165 6.655 91.425 ;
        RECT 6.735 91.165 6.995 91.425 ;
        RECT 7.055 91.165 7.315 91.425 ;
        RECT 7.460 91.165 7.720 91.425 ;
        RECT 7.800 91.165 8.060 91.425 ;
        RECT 8.250 91.165 8.510 91.425 ;
        RECT 8.590 91.165 8.850 91.425 ;
        RECT 8.910 91.165 9.170 91.425 ;
        RECT 9.315 91.165 9.575 91.425 ;
        RECT 9.655 91.165 9.915 91.425 ;
        RECT 62.945 91.360 63.205 91.620 ;
        RECT 63.285 91.360 63.545 91.620 ;
        RECT 63.850 91.360 64.110 91.620 ;
        RECT 64.190 91.360 64.450 91.620 ;
        RECT 64.510 91.360 64.770 91.620 ;
        RECT 64.915 91.360 65.175 91.620 ;
        RECT 65.255 91.360 65.515 91.620 ;
        RECT 65.575 91.360 65.835 91.620 ;
        RECT 66.060 91.360 66.320 91.620 ;
        RECT 4.660 80.725 4.920 80.985 ;
        RECT 5.000 80.725 5.260 80.985 ;
        RECT 5.320 80.725 5.580 80.985 ;
        RECT 5.725 80.725 5.985 80.985 ;
        RECT 6.065 80.725 6.325 80.985 ;
        RECT 6.385 80.725 6.645 80.985 ;
        RECT 6.870 80.725 7.130 80.985 ;
        RECT 7.210 80.725 7.470 80.985 ;
        RECT 7.530 80.725 7.790 80.985 ;
        RECT 7.935 80.725 8.195 80.985 ;
        RECT 8.275 80.725 8.535 80.985 ;
        RECT 4.660 80.400 4.920 80.660 ;
        RECT 5.000 80.400 5.260 80.660 ;
        RECT 5.320 80.400 5.580 80.660 ;
        RECT 5.725 80.400 5.985 80.660 ;
        RECT 6.065 80.400 6.325 80.660 ;
        RECT 6.385 80.400 6.645 80.660 ;
        RECT 6.870 80.400 7.130 80.660 ;
        RECT 7.210 80.400 7.470 80.660 ;
        RECT 7.530 80.400 7.790 80.660 ;
        RECT 7.935 80.400 8.195 80.660 ;
        RECT 8.275 80.400 8.535 80.660 ;
        RECT 4.660 80.070 4.920 80.330 ;
        RECT 5.000 80.070 5.260 80.330 ;
        RECT 5.320 80.070 5.580 80.330 ;
        RECT 5.725 80.070 5.985 80.330 ;
        RECT 6.065 80.070 6.325 80.330 ;
        RECT 6.385 80.070 6.645 80.330 ;
        RECT 6.870 80.070 7.130 80.330 ;
        RECT 7.210 80.070 7.470 80.330 ;
        RECT 7.530 80.070 7.790 80.330 ;
        RECT 7.935 80.070 8.195 80.330 ;
        RECT 8.275 80.070 8.535 80.330 ;
        RECT 4.660 79.670 4.920 79.930 ;
        RECT 5.000 79.670 5.260 79.930 ;
        RECT 5.320 79.670 5.580 79.930 ;
        RECT 5.725 79.670 5.985 79.930 ;
        RECT 6.065 79.670 6.325 79.930 ;
        RECT 6.385 79.670 6.645 79.930 ;
        RECT 6.870 79.670 7.130 79.930 ;
        RECT 7.210 79.670 7.470 79.930 ;
        RECT 7.530 79.670 7.790 79.930 ;
        RECT 7.935 79.670 8.195 79.930 ;
        RECT 8.275 79.670 8.535 79.930 ;
        RECT 4.660 79.345 4.920 79.605 ;
        RECT 5.000 79.345 5.260 79.605 ;
        RECT 5.320 79.345 5.580 79.605 ;
        RECT 5.725 79.345 5.985 79.605 ;
        RECT 6.065 79.345 6.325 79.605 ;
        RECT 6.385 79.345 6.645 79.605 ;
        RECT 6.870 79.345 7.130 79.605 ;
        RECT 7.210 79.345 7.470 79.605 ;
        RECT 7.530 79.345 7.790 79.605 ;
        RECT 7.935 79.345 8.195 79.605 ;
        RECT 8.275 79.345 8.535 79.605 ;
        RECT 4.660 79.015 4.920 79.275 ;
        RECT 5.000 79.015 5.260 79.275 ;
        RECT 5.320 79.015 5.580 79.275 ;
        RECT 5.725 79.015 5.985 79.275 ;
        RECT 6.065 79.015 6.325 79.275 ;
        RECT 6.385 79.015 6.645 79.275 ;
        RECT 6.870 79.015 7.130 79.275 ;
        RECT 7.210 79.015 7.470 79.275 ;
        RECT 7.530 79.015 7.790 79.275 ;
        RECT 7.935 79.015 8.195 79.275 ;
        RECT 8.275 79.015 8.535 79.275 ;
        RECT 4.660 78.545 4.920 78.805 ;
        RECT 5.000 78.545 5.260 78.805 ;
        RECT 5.320 78.545 5.580 78.805 ;
        RECT 5.725 78.545 5.985 78.805 ;
        RECT 6.065 78.545 6.325 78.805 ;
        RECT 6.385 78.545 6.645 78.805 ;
        RECT 6.870 78.545 7.130 78.805 ;
        RECT 7.210 78.545 7.470 78.805 ;
        RECT 7.530 78.545 7.790 78.805 ;
        RECT 7.935 78.545 8.195 78.805 ;
        RECT 8.275 78.545 8.535 78.805 ;
        RECT 4.660 78.220 4.920 78.480 ;
        RECT 5.000 78.220 5.260 78.480 ;
        RECT 5.320 78.220 5.580 78.480 ;
        RECT 5.725 78.220 5.985 78.480 ;
        RECT 6.065 78.220 6.325 78.480 ;
        RECT 6.385 78.220 6.645 78.480 ;
        RECT 6.870 78.220 7.130 78.480 ;
        RECT 7.210 78.220 7.470 78.480 ;
        RECT 7.530 78.220 7.790 78.480 ;
        RECT 7.935 78.220 8.195 78.480 ;
        RECT 8.275 78.220 8.535 78.480 ;
        RECT 4.660 77.890 4.920 78.150 ;
        RECT 5.000 77.890 5.260 78.150 ;
        RECT 5.320 77.890 5.580 78.150 ;
        RECT 5.725 77.890 5.985 78.150 ;
        RECT 6.065 77.890 6.325 78.150 ;
        RECT 6.385 77.890 6.645 78.150 ;
        RECT 6.870 77.890 7.130 78.150 ;
        RECT 7.210 77.890 7.470 78.150 ;
        RECT 7.530 77.890 7.790 78.150 ;
        RECT 7.935 77.890 8.195 78.150 ;
        RECT 8.275 77.890 8.535 78.150 ;
        RECT 4.660 77.490 4.920 77.750 ;
        RECT 5.000 77.490 5.260 77.750 ;
        RECT 5.320 77.490 5.580 77.750 ;
        RECT 5.725 77.490 5.985 77.750 ;
        RECT 6.065 77.490 6.325 77.750 ;
        RECT 6.385 77.490 6.645 77.750 ;
        RECT 6.870 77.490 7.130 77.750 ;
        RECT 7.210 77.490 7.470 77.750 ;
        RECT 7.530 77.490 7.790 77.750 ;
        RECT 7.935 77.490 8.195 77.750 ;
        RECT 8.275 77.490 8.535 77.750 ;
        RECT 4.660 77.165 4.920 77.425 ;
        RECT 5.000 77.165 5.260 77.425 ;
        RECT 5.320 77.165 5.580 77.425 ;
        RECT 5.725 77.165 5.985 77.425 ;
        RECT 6.065 77.165 6.325 77.425 ;
        RECT 6.385 77.165 6.645 77.425 ;
        RECT 6.870 77.165 7.130 77.425 ;
        RECT 7.210 77.165 7.470 77.425 ;
        RECT 7.530 77.165 7.790 77.425 ;
        RECT 7.935 77.165 8.195 77.425 ;
        RECT 8.275 77.165 8.535 77.425 ;
        RECT 62.130 77.215 62.390 77.475 ;
        RECT 62.470 77.215 62.730 77.475 ;
        RECT 63.035 77.215 63.295 77.475 ;
        RECT 63.375 77.215 63.635 77.475 ;
        RECT 63.695 77.215 63.955 77.475 ;
        RECT 64.100 77.215 64.360 77.475 ;
        RECT 64.440 77.215 64.700 77.475 ;
        RECT 64.760 77.215 65.020 77.475 ;
        RECT 65.245 77.215 65.505 77.475 ;
        RECT 65.865 77.215 66.125 77.475 ;
        RECT 66.205 77.215 66.465 77.475 ;
        RECT 66.525 77.215 66.785 77.475 ;
        RECT 67.010 77.215 67.270 77.475 ;
        RECT 4.660 76.835 4.920 77.095 ;
        RECT 5.000 76.835 5.260 77.095 ;
        RECT 5.320 76.835 5.580 77.095 ;
        RECT 5.725 76.835 5.985 77.095 ;
        RECT 6.065 76.835 6.325 77.095 ;
        RECT 6.385 76.835 6.645 77.095 ;
        RECT 6.870 76.835 7.130 77.095 ;
        RECT 7.210 76.835 7.470 77.095 ;
        RECT 7.530 76.835 7.790 77.095 ;
        RECT 7.935 76.835 8.195 77.095 ;
        RECT 8.275 76.835 8.535 77.095 ;
        RECT 62.130 76.890 62.390 77.150 ;
        RECT 62.470 76.890 62.730 77.150 ;
        RECT 63.035 76.890 63.295 77.150 ;
        RECT 63.375 76.890 63.635 77.150 ;
        RECT 63.695 76.890 63.955 77.150 ;
        RECT 64.100 76.890 64.360 77.150 ;
        RECT 64.440 76.890 64.700 77.150 ;
        RECT 64.760 76.890 65.020 77.150 ;
        RECT 65.245 76.890 65.505 77.150 ;
        RECT 65.865 76.890 66.125 77.150 ;
        RECT 66.205 76.890 66.465 77.150 ;
        RECT 66.525 76.890 66.785 77.150 ;
        RECT 67.010 76.890 67.270 77.150 ;
        RECT 4.660 76.305 4.920 76.565 ;
        RECT 5.000 76.305 5.260 76.565 ;
        RECT 5.320 76.305 5.580 76.565 ;
        RECT 5.725 76.305 5.985 76.565 ;
        RECT 6.065 76.305 6.325 76.565 ;
        RECT 6.385 76.305 6.645 76.565 ;
        RECT 6.870 76.305 7.130 76.565 ;
        RECT 7.210 76.305 7.470 76.565 ;
        RECT 7.530 76.305 7.790 76.565 ;
        RECT 7.935 76.305 8.195 76.565 ;
        RECT 8.275 76.305 8.535 76.565 ;
        RECT 62.130 76.465 62.390 76.725 ;
        RECT 62.470 76.465 62.730 76.725 ;
        RECT 63.035 76.465 63.295 76.725 ;
        RECT 63.375 76.465 63.635 76.725 ;
        RECT 63.695 76.465 63.955 76.725 ;
        RECT 64.100 76.465 64.360 76.725 ;
        RECT 64.440 76.465 64.700 76.725 ;
        RECT 64.760 76.465 65.020 76.725 ;
        RECT 65.245 76.465 65.505 76.725 ;
        RECT 65.865 76.465 66.125 76.725 ;
        RECT 66.205 76.465 66.465 76.725 ;
        RECT 66.525 76.465 66.785 76.725 ;
        RECT 67.010 76.465 67.270 76.725 ;
        RECT 4.660 75.980 4.920 76.240 ;
        RECT 5.000 75.980 5.260 76.240 ;
        RECT 5.320 75.980 5.580 76.240 ;
        RECT 5.725 75.980 5.985 76.240 ;
        RECT 6.065 75.980 6.325 76.240 ;
        RECT 6.385 75.980 6.645 76.240 ;
        RECT 6.870 75.980 7.130 76.240 ;
        RECT 7.210 75.980 7.470 76.240 ;
        RECT 7.530 75.980 7.790 76.240 ;
        RECT 7.935 75.980 8.195 76.240 ;
        RECT 8.275 75.980 8.535 76.240 ;
        RECT 62.130 76.140 62.390 76.400 ;
        RECT 62.470 76.140 62.730 76.400 ;
        RECT 63.035 76.140 63.295 76.400 ;
        RECT 63.375 76.140 63.635 76.400 ;
        RECT 63.695 76.140 63.955 76.400 ;
        RECT 64.100 76.140 64.360 76.400 ;
        RECT 64.440 76.140 64.700 76.400 ;
        RECT 64.760 76.140 65.020 76.400 ;
        RECT 65.245 76.140 65.505 76.400 ;
        RECT 65.865 76.140 66.125 76.400 ;
        RECT 66.205 76.140 66.465 76.400 ;
        RECT 66.525 76.140 66.785 76.400 ;
        RECT 67.010 76.140 67.270 76.400 ;
        RECT 4.660 75.650 4.920 75.910 ;
        RECT 5.000 75.650 5.260 75.910 ;
        RECT 5.320 75.650 5.580 75.910 ;
        RECT 5.725 75.650 5.985 75.910 ;
        RECT 6.065 75.650 6.325 75.910 ;
        RECT 6.385 75.650 6.645 75.910 ;
        RECT 6.870 75.650 7.130 75.910 ;
        RECT 7.210 75.650 7.470 75.910 ;
        RECT 7.530 75.650 7.790 75.910 ;
        RECT 7.935 75.650 8.195 75.910 ;
        RECT 8.275 75.650 8.535 75.910 ;
        RECT 62.130 75.715 62.390 75.975 ;
        RECT 62.470 75.715 62.730 75.975 ;
        RECT 63.035 75.715 63.295 75.975 ;
        RECT 63.375 75.715 63.635 75.975 ;
        RECT 63.695 75.715 63.955 75.975 ;
        RECT 64.100 75.715 64.360 75.975 ;
        RECT 64.440 75.715 64.700 75.975 ;
        RECT 64.760 75.715 65.020 75.975 ;
        RECT 65.245 75.715 65.505 75.975 ;
        RECT 65.865 75.715 66.125 75.975 ;
        RECT 66.205 75.715 66.465 75.975 ;
        RECT 66.525 75.715 66.785 75.975 ;
        RECT 67.010 75.715 67.270 75.975 ;
        RECT 4.660 75.250 4.920 75.510 ;
        RECT 5.000 75.250 5.260 75.510 ;
        RECT 5.320 75.250 5.580 75.510 ;
        RECT 5.725 75.250 5.985 75.510 ;
        RECT 6.065 75.250 6.325 75.510 ;
        RECT 6.385 75.250 6.645 75.510 ;
        RECT 6.870 75.250 7.130 75.510 ;
        RECT 7.210 75.250 7.470 75.510 ;
        RECT 7.530 75.250 7.790 75.510 ;
        RECT 7.935 75.250 8.195 75.510 ;
        RECT 8.275 75.250 8.535 75.510 ;
        RECT 62.130 75.390 62.390 75.650 ;
        RECT 62.470 75.390 62.730 75.650 ;
        RECT 63.035 75.390 63.295 75.650 ;
        RECT 63.375 75.390 63.635 75.650 ;
        RECT 63.695 75.390 63.955 75.650 ;
        RECT 64.100 75.390 64.360 75.650 ;
        RECT 64.440 75.390 64.700 75.650 ;
        RECT 64.760 75.390 65.020 75.650 ;
        RECT 65.245 75.390 65.505 75.650 ;
        RECT 65.865 75.390 66.125 75.650 ;
        RECT 66.205 75.390 66.465 75.650 ;
        RECT 66.525 75.390 66.785 75.650 ;
        RECT 67.010 75.390 67.270 75.650 ;
        RECT 4.660 74.925 4.920 75.185 ;
        RECT 5.000 74.925 5.260 75.185 ;
        RECT 5.320 74.925 5.580 75.185 ;
        RECT 5.725 74.925 5.985 75.185 ;
        RECT 6.065 74.925 6.325 75.185 ;
        RECT 6.385 74.925 6.645 75.185 ;
        RECT 6.870 74.925 7.130 75.185 ;
        RECT 7.210 74.925 7.470 75.185 ;
        RECT 7.530 74.925 7.790 75.185 ;
        RECT 7.935 74.925 8.195 75.185 ;
        RECT 8.275 74.925 8.535 75.185 ;
        RECT 62.130 74.925 62.390 75.185 ;
        RECT 62.470 74.925 62.730 75.185 ;
        RECT 63.035 74.925 63.295 75.185 ;
        RECT 63.375 74.925 63.635 75.185 ;
        RECT 63.695 74.925 63.955 75.185 ;
        RECT 64.100 74.925 64.360 75.185 ;
        RECT 64.440 74.925 64.700 75.185 ;
        RECT 64.760 74.925 65.020 75.185 ;
        RECT 65.245 74.925 65.505 75.185 ;
        RECT 65.865 74.925 66.125 75.185 ;
        RECT 66.205 74.925 66.465 75.185 ;
        RECT 66.525 74.925 66.785 75.185 ;
        RECT 67.010 74.925 67.270 75.185 ;
        RECT 4.660 74.595 4.920 74.855 ;
        RECT 5.000 74.595 5.260 74.855 ;
        RECT 5.320 74.595 5.580 74.855 ;
        RECT 5.725 74.595 5.985 74.855 ;
        RECT 6.065 74.595 6.325 74.855 ;
        RECT 6.385 74.595 6.645 74.855 ;
        RECT 6.870 74.595 7.130 74.855 ;
        RECT 7.210 74.595 7.470 74.855 ;
        RECT 7.530 74.595 7.790 74.855 ;
        RECT 7.935 74.595 8.195 74.855 ;
        RECT 8.275 74.595 8.535 74.855 ;
        RECT 62.130 74.600 62.390 74.860 ;
        RECT 62.470 74.600 62.730 74.860 ;
        RECT 63.035 74.600 63.295 74.860 ;
        RECT 63.375 74.600 63.635 74.860 ;
        RECT 63.695 74.600 63.955 74.860 ;
        RECT 64.100 74.600 64.360 74.860 ;
        RECT 64.440 74.600 64.700 74.860 ;
        RECT 64.760 74.600 65.020 74.860 ;
        RECT 65.245 74.600 65.505 74.860 ;
        RECT 65.865 74.600 66.125 74.860 ;
        RECT 66.205 74.600 66.465 74.860 ;
        RECT 66.525 74.600 66.785 74.860 ;
        RECT 67.010 74.600 67.270 74.860 ;
        RECT 4.660 74.125 4.920 74.385 ;
        RECT 5.000 74.125 5.260 74.385 ;
        RECT 5.320 74.125 5.580 74.385 ;
        RECT 5.725 74.125 5.985 74.385 ;
        RECT 6.065 74.125 6.325 74.385 ;
        RECT 6.385 74.125 6.645 74.385 ;
        RECT 6.870 74.125 7.130 74.385 ;
        RECT 7.210 74.125 7.470 74.385 ;
        RECT 7.530 74.125 7.790 74.385 ;
        RECT 7.935 74.125 8.195 74.385 ;
        RECT 8.275 74.125 8.535 74.385 ;
        RECT 4.660 73.800 4.920 74.060 ;
        RECT 5.000 73.800 5.260 74.060 ;
        RECT 5.320 73.800 5.580 74.060 ;
        RECT 5.725 73.800 5.985 74.060 ;
        RECT 6.065 73.800 6.325 74.060 ;
        RECT 6.385 73.800 6.645 74.060 ;
        RECT 6.870 73.800 7.130 74.060 ;
        RECT 7.210 73.800 7.470 74.060 ;
        RECT 7.530 73.800 7.790 74.060 ;
        RECT 7.935 73.800 8.195 74.060 ;
        RECT 8.275 73.800 8.535 74.060 ;
        RECT 4.660 73.470 4.920 73.730 ;
        RECT 5.000 73.470 5.260 73.730 ;
        RECT 5.320 73.470 5.580 73.730 ;
        RECT 5.725 73.470 5.985 73.730 ;
        RECT 6.065 73.470 6.325 73.730 ;
        RECT 6.385 73.470 6.645 73.730 ;
        RECT 6.870 73.470 7.130 73.730 ;
        RECT 7.210 73.470 7.470 73.730 ;
        RECT 7.530 73.470 7.790 73.730 ;
        RECT 7.935 73.470 8.195 73.730 ;
        RECT 8.275 73.470 8.535 73.730 ;
        RECT 4.660 73.070 4.920 73.330 ;
        RECT 5.000 73.070 5.260 73.330 ;
        RECT 5.320 73.070 5.580 73.330 ;
        RECT 5.725 73.070 5.985 73.330 ;
        RECT 6.065 73.070 6.325 73.330 ;
        RECT 6.385 73.070 6.645 73.330 ;
        RECT 6.870 73.070 7.130 73.330 ;
        RECT 7.210 73.070 7.470 73.330 ;
        RECT 7.530 73.070 7.790 73.330 ;
        RECT 7.935 73.070 8.195 73.330 ;
        RECT 8.275 73.070 8.535 73.330 ;
      LAYER met2 ;
        RECT 4.160 157.300 17.700 165.310 ;
        RECT 4.160 72.730 11.050 157.300 ;
        RECT 62.700 112.325 67.900 114.325 ;
        RECT 62.700 93.125 64.700 112.325 ;
        RECT 62.275 90.875 66.710 93.125 ;
        RECT 62.700 77.705 64.700 90.875 ;
        RECT 61.810 74.405 67.560 77.705 ;
    END
  END vssio
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 14.880 38.600 15.310 39.385 ;
        RECT 25.460 38.600 25.890 39.385 ;
        RECT 44.320 38.600 44.750 39.385 ;
        RECT 63.180 38.600 63.610 39.385 ;
        RECT 12.805 28.255 13.235 29.040 ;
        RECT 29.365 28.255 29.795 29.040 ;
        RECT 39.945 28.255 40.375 29.040 ;
        RECT 54.205 28.255 54.635 29.040 ;
        RECT 55.390 27.700 73.060 29.070 ;
        RECT 55.190 27.270 73.210 27.700 ;
      LAYER li1 ;
        RECT 14.950 38.495 15.240 39.220 ;
        RECT 17.860 38.495 18.030 38.955 ;
        RECT 18.700 38.495 18.870 38.955 ;
        RECT 21.435 38.495 21.700 38.955 ;
        RECT 22.370 38.495 22.540 38.955 ;
        RECT 23.210 38.495 23.460 38.960 ;
        RECT 25.530 38.495 25.820 39.220 ;
        RECT 27.890 38.495 28.140 38.960 ;
        RECT 28.810 38.495 28.980 38.955 ;
        RECT 29.650 38.495 29.915 38.955 ;
        RECT 32.480 38.495 32.650 38.955 ;
        RECT 33.320 38.495 33.490 38.955 ;
        RECT 36.170 38.495 36.420 38.960 ;
        RECT 37.090 38.495 37.260 38.955 ;
        RECT 37.930 38.495 38.195 38.955 ;
        RECT 42.700 38.495 42.870 38.955 ;
        RECT 43.540 38.495 43.710 38.955 ;
        RECT 44.390 38.495 44.680 39.220 ;
        RECT 46.750 38.495 47.000 38.960 ;
        RECT 47.670 38.495 47.840 38.955 ;
        RECT 48.510 38.495 48.775 38.955 ;
        RECT 51.340 38.495 51.510 38.955 ;
        RECT 52.180 38.495 52.350 38.955 ;
        RECT 55.030 38.495 55.280 38.960 ;
        RECT 55.950 38.495 56.120 38.955 ;
        RECT 56.790 38.495 57.055 38.955 ;
        RECT 59.620 38.495 59.790 38.955 ;
        RECT 60.460 38.495 60.630 38.955 ;
        RECT 63.250 38.495 63.540 39.220 ;
        RECT 14.865 38.325 63.625 38.495 ;
        RECT 12.875 28.150 13.165 28.875 ;
        RECT 15.235 28.150 15.485 28.615 ;
        RECT 16.155 28.150 16.325 28.610 ;
        RECT 16.995 28.150 17.260 28.610 ;
        RECT 19.530 28.150 19.815 28.620 ;
        RECT 20.485 28.150 20.655 28.620 ;
        RECT 21.325 28.150 21.495 28.620 ;
        RECT 22.165 28.150 22.335 28.620 ;
        RECT 23.005 28.150 23.280 28.970 ;
        RECT 25.355 28.150 25.605 28.615 ;
        RECT 26.275 28.150 26.445 28.610 ;
        RECT 27.115 28.150 27.380 28.610 ;
        RECT 29.435 28.150 29.725 28.875 ;
        RECT 31.795 28.150 32.045 28.615 ;
        RECT 32.715 28.150 32.885 28.610 ;
        RECT 33.555 28.150 33.820 28.610 ;
        RECT 36.090 28.150 36.375 28.620 ;
        RECT 37.045 28.150 37.215 28.620 ;
        RECT 37.885 28.150 38.055 28.620 ;
        RECT 38.725 28.150 38.895 28.620 ;
        RECT 39.565 28.150 39.840 28.970 ;
        RECT 40.015 28.150 40.305 28.875 ;
        RECT 46.055 28.150 46.305 28.615 ;
        RECT 46.975 28.150 47.145 28.610 ;
        RECT 47.815 28.150 48.080 28.610 ;
        RECT 50.350 28.150 50.635 28.620 ;
        RECT 51.305 28.150 51.475 28.620 ;
        RECT 52.145 28.150 52.315 28.620 ;
        RECT 52.985 28.150 53.155 28.620 ;
        RECT 53.825 28.150 54.100 28.970 ;
        RECT 54.275 28.150 54.565 28.875 ;
        RECT 12.790 27.980 54.650 28.150 ;
        RECT 55.480 27.910 56.010 28.980 ;
        RECT 56.760 27.910 57.650 28.880 ;
        RECT 58.320 27.910 59.210 28.880 ;
        RECT 59.880 27.910 60.770 28.880 ;
        RECT 61.440 27.910 62.330 28.880 ;
        RECT 63.000 27.910 63.890 28.880 ;
        RECT 64.560 27.910 65.450 28.880 ;
        RECT 66.120 27.910 67.010 28.880 ;
        RECT 67.750 27.910 68.640 28.510 ;
        RECT 69.225 27.910 70.120 28.510 ;
        RECT 70.850 27.900 71.740 28.510 ;
        RECT 72.435 27.910 72.970 28.895 ;
        RECT 55.320 27.400 73.080 27.570 ;
      LAYER mcon ;
        RECT 15.010 38.325 15.180 38.495 ;
        RECT 15.470 38.325 15.640 38.495 ;
        RECT 15.930 38.325 16.100 38.495 ;
        RECT 16.390 38.325 16.560 38.495 ;
        RECT 16.850 38.325 17.020 38.495 ;
        RECT 17.310 38.325 17.480 38.495 ;
        RECT 17.770 38.325 17.940 38.495 ;
        RECT 18.230 38.325 18.400 38.495 ;
        RECT 18.690 38.325 18.860 38.495 ;
        RECT 19.150 38.325 19.320 38.495 ;
        RECT 19.610 38.325 19.780 38.495 ;
        RECT 20.070 38.325 20.240 38.495 ;
        RECT 20.530 38.325 20.700 38.495 ;
        RECT 20.990 38.325 21.160 38.495 ;
        RECT 21.450 38.325 21.620 38.495 ;
        RECT 21.910 38.325 22.080 38.495 ;
        RECT 22.370 38.325 22.540 38.495 ;
        RECT 22.830 38.325 23.000 38.495 ;
        RECT 23.290 38.325 23.460 38.495 ;
        RECT 23.750 38.325 23.920 38.495 ;
        RECT 24.210 38.325 24.380 38.495 ;
        RECT 24.670 38.325 24.840 38.495 ;
        RECT 25.130 38.325 25.300 38.495 ;
        RECT 25.590 38.325 25.760 38.495 ;
        RECT 26.050 38.325 26.220 38.495 ;
        RECT 26.510 38.325 26.680 38.495 ;
        RECT 26.970 38.325 27.140 38.495 ;
        RECT 27.430 38.325 27.600 38.495 ;
        RECT 27.890 38.325 28.060 38.495 ;
        RECT 28.350 38.325 28.520 38.495 ;
        RECT 28.810 38.325 28.980 38.495 ;
        RECT 29.270 38.325 29.440 38.495 ;
        RECT 29.730 38.325 29.900 38.495 ;
        RECT 30.190 38.325 30.360 38.495 ;
        RECT 30.650 38.325 30.820 38.495 ;
        RECT 31.110 38.325 31.280 38.495 ;
        RECT 31.570 38.325 31.740 38.495 ;
        RECT 32.030 38.325 32.200 38.495 ;
        RECT 32.490 38.325 32.660 38.495 ;
        RECT 32.950 38.325 33.120 38.495 ;
        RECT 33.410 38.325 33.580 38.495 ;
        RECT 33.870 38.325 34.040 38.495 ;
        RECT 34.330 38.325 34.500 38.495 ;
        RECT 34.790 38.325 34.960 38.495 ;
        RECT 35.250 38.325 35.420 38.495 ;
        RECT 35.710 38.325 35.880 38.495 ;
        RECT 36.170 38.325 36.340 38.495 ;
        RECT 36.630 38.325 36.800 38.495 ;
        RECT 37.090 38.325 37.260 38.495 ;
        RECT 37.550 38.325 37.720 38.495 ;
        RECT 38.010 38.325 38.180 38.495 ;
        RECT 38.470 38.325 38.640 38.495 ;
        RECT 38.930 38.325 39.100 38.495 ;
        RECT 39.390 38.325 39.560 38.495 ;
        RECT 39.850 38.325 40.020 38.495 ;
        RECT 40.310 38.325 40.480 38.495 ;
        RECT 40.770 38.325 40.940 38.495 ;
        RECT 41.230 38.325 41.400 38.495 ;
        RECT 41.690 38.325 41.860 38.495 ;
        RECT 42.150 38.325 42.320 38.495 ;
        RECT 42.610 38.325 42.780 38.495 ;
        RECT 43.070 38.325 43.240 38.495 ;
        RECT 43.530 38.325 43.700 38.495 ;
        RECT 43.990 38.325 44.160 38.495 ;
        RECT 44.450 38.325 44.620 38.495 ;
        RECT 44.910 38.325 45.080 38.495 ;
        RECT 45.370 38.325 45.540 38.495 ;
        RECT 45.830 38.325 46.000 38.495 ;
        RECT 46.290 38.325 46.460 38.495 ;
        RECT 46.750 38.325 46.920 38.495 ;
        RECT 47.210 38.325 47.380 38.495 ;
        RECT 47.670 38.325 47.840 38.495 ;
        RECT 48.130 38.325 48.300 38.495 ;
        RECT 48.590 38.325 48.760 38.495 ;
        RECT 49.050 38.325 49.220 38.495 ;
        RECT 49.510 38.325 49.680 38.495 ;
        RECT 49.970 38.325 50.140 38.495 ;
        RECT 50.430 38.325 50.600 38.495 ;
        RECT 50.890 38.325 51.060 38.495 ;
        RECT 51.350 38.325 51.520 38.495 ;
        RECT 51.810 38.325 51.980 38.495 ;
        RECT 52.270 38.325 52.440 38.495 ;
        RECT 52.730 38.325 52.900 38.495 ;
        RECT 53.190 38.325 53.360 38.495 ;
        RECT 53.650 38.325 53.820 38.495 ;
        RECT 54.110 38.325 54.280 38.495 ;
        RECT 54.570 38.325 54.740 38.495 ;
        RECT 55.030 38.325 55.200 38.495 ;
        RECT 55.490 38.325 55.660 38.495 ;
        RECT 55.950 38.325 56.120 38.495 ;
        RECT 56.410 38.325 56.580 38.495 ;
        RECT 56.870 38.325 57.040 38.495 ;
        RECT 57.330 38.325 57.500 38.495 ;
        RECT 57.790 38.325 57.960 38.495 ;
        RECT 58.250 38.325 58.420 38.495 ;
        RECT 58.710 38.325 58.880 38.495 ;
        RECT 59.170 38.325 59.340 38.495 ;
        RECT 59.630 38.325 59.800 38.495 ;
        RECT 60.090 38.325 60.260 38.495 ;
        RECT 60.550 38.325 60.720 38.495 ;
        RECT 61.010 38.325 61.180 38.495 ;
        RECT 61.470 38.325 61.640 38.495 ;
        RECT 61.930 38.325 62.100 38.495 ;
        RECT 62.390 38.325 62.560 38.495 ;
        RECT 62.850 38.325 63.020 38.495 ;
        RECT 63.310 38.325 63.480 38.495 ;
        RECT 12.935 27.980 13.105 28.150 ;
        RECT 13.395 27.980 13.565 28.150 ;
        RECT 13.855 27.980 14.025 28.150 ;
        RECT 14.315 27.980 14.485 28.150 ;
        RECT 14.775 27.980 14.945 28.150 ;
        RECT 15.235 27.980 15.405 28.150 ;
        RECT 15.695 27.980 15.865 28.150 ;
        RECT 16.155 27.980 16.325 28.150 ;
        RECT 16.615 27.980 16.785 28.150 ;
        RECT 17.075 27.980 17.245 28.150 ;
        RECT 17.535 27.980 17.705 28.150 ;
        RECT 17.995 27.980 18.165 28.150 ;
        RECT 18.455 27.980 18.625 28.150 ;
        RECT 18.915 27.980 19.085 28.150 ;
        RECT 19.375 27.980 19.545 28.150 ;
        RECT 19.835 27.980 20.005 28.150 ;
        RECT 20.295 27.980 20.465 28.150 ;
        RECT 20.755 27.980 20.925 28.150 ;
        RECT 21.215 27.980 21.385 28.150 ;
        RECT 21.675 27.980 21.845 28.150 ;
        RECT 22.135 27.980 22.305 28.150 ;
        RECT 22.595 27.980 22.765 28.150 ;
        RECT 23.055 27.980 23.225 28.150 ;
        RECT 23.515 27.980 23.685 28.150 ;
        RECT 23.975 27.980 24.145 28.150 ;
        RECT 24.435 27.980 24.605 28.150 ;
        RECT 24.895 27.980 25.065 28.150 ;
        RECT 25.355 27.980 25.525 28.150 ;
        RECT 25.815 27.980 25.985 28.150 ;
        RECT 26.275 27.980 26.445 28.150 ;
        RECT 26.735 27.980 26.905 28.150 ;
        RECT 27.195 27.980 27.365 28.150 ;
        RECT 27.655 27.980 27.825 28.150 ;
        RECT 28.115 27.980 28.285 28.150 ;
        RECT 28.575 27.980 28.745 28.150 ;
        RECT 29.035 27.980 29.205 28.150 ;
        RECT 29.495 27.980 29.665 28.150 ;
        RECT 29.955 27.980 30.125 28.150 ;
        RECT 30.415 27.980 30.585 28.150 ;
        RECT 30.875 27.980 31.045 28.150 ;
        RECT 31.335 27.980 31.505 28.150 ;
        RECT 31.795 27.980 31.965 28.150 ;
        RECT 32.255 27.980 32.425 28.150 ;
        RECT 32.715 27.980 32.885 28.150 ;
        RECT 33.175 27.980 33.345 28.150 ;
        RECT 33.635 27.980 33.805 28.150 ;
        RECT 34.095 27.980 34.265 28.150 ;
        RECT 34.555 27.980 34.725 28.150 ;
        RECT 35.015 27.980 35.185 28.150 ;
        RECT 35.475 27.980 35.645 28.150 ;
        RECT 35.935 27.980 36.105 28.150 ;
        RECT 36.395 27.980 36.565 28.150 ;
        RECT 36.855 27.980 37.025 28.150 ;
        RECT 37.315 27.980 37.485 28.150 ;
        RECT 37.775 27.980 37.945 28.150 ;
        RECT 38.235 27.980 38.405 28.150 ;
        RECT 38.695 27.980 38.865 28.150 ;
        RECT 39.155 27.980 39.325 28.150 ;
        RECT 39.615 27.980 39.785 28.150 ;
        RECT 40.075 27.980 40.245 28.150 ;
        RECT 40.535 27.980 40.705 28.150 ;
        RECT 40.995 27.980 41.165 28.150 ;
        RECT 41.455 27.980 41.625 28.150 ;
        RECT 41.915 27.980 42.085 28.150 ;
        RECT 42.375 27.980 42.545 28.150 ;
        RECT 42.835 27.980 43.005 28.150 ;
        RECT 43.295 27.980 43.465 28.150 ;
        RECT 43.755 27.980 43.925 28.150 ;
        RECT 44.215 27.980 44.385 28.150 ;
        RECT 44.675 27.980 44.845 28.150 ;
        RECT 45.135 27.980 45.305 28.150 ;
        RECT 45.595 27.980 45.765 28.150 ;
        RECT 46.055 27.980 46.225 28.150 ;
        RECT 46.515 27.980 46.685 28.150 ;
        RECT 46.975 27.980 47.145 28.150 ;
        RECT 47.435 27.980 47.605 28.150 ;
        RECT 47.895 27.980 48.065 28.150 ;
        RECT 48.355 27.980 48.525 28.150 ;
        RECT 48.815 27.980 48.985 28.150 ;
        RECT 49.275 27.980 49.445 28.150 ;
        RECT 49.735 27.980 49.905 28.150 ;
        RECT 50.195 27.980 50.365 28.150 ;
        RECT 50.655 27.980 50.825 28.150 ;
        RECT 51.115 27.980 51.285 28.150 ;
        RECT 51.575 27.980 51.745 28.150 ;
        RECT 52.035 27.980 52.205 28.150 ;
        RECT 52.495 27.980 52.665 28.150 ;
        RECT 52.955 27.980 53.125 28.150 ;
        RECT 53.415 27.980 53.585 28.150 ;
        RECT 53.875 27.980 54.045 28.150 ;
        RECT 54.335 27.980 54.505 28.150 ;
        RECT 55.840 27.910 56.010 28.080 ;
        RECT 57.120 27.910 57.290 28.080 ;
        RECT 57.480 27.910 57.650 28.080 ;
        RECT 58.680 27.910 58.850 28.080 ;
        RECT 59.040 27.910 59.210 28.080 ;
        RECT 60.240 27.910 60.410 28.080 ;
        RECT 60.600 27.910 60.770 28.080 ;
        RECT 61.800 27.910 61.970 28.080 ;
        RECT 62.160 27.910 62.330 28.080 ;
        RECT 63.360 27.910 63.530 28.080 ;
        RECT 63.720 27.910 63.890 28.080 ;
        RECT 64.920 27.910 65.090 28.080 ;
        RECT 65.280 27.910 65.450 28.080 ;
        RECT 66.480 27.910 66.650 28.080 ;
        RECT 66.840 27.910 67.010 28.080 ;
        RECT 68.110 27.910 68.280 28.080 ;
        RECT 68.470 27.910 68.640 28.080 ;
        RECT 69.230 27.910 69.400 28.080 ;
        RECT 69.590 27.910 69.760 28.080 ;
        RECT 69.950 27.910 70.120 28.080 ;
        RECT 70.850 27.910 71.020 28.080 ;
        RECT 71.210 27.910 71.380 28.080 ;
        RECT 71.570 27.910 71.740 28.080 ;
        RECT 72.795 27.910 72.965 28.080 ;
        RECT 55.475 27.400 55.645 27.570 ;
        RECT 55.955 27.400 56.125 27.570 ;
        RECT 56.435 27.400 56.605 27.570 ;
        RECT 56.915 27.400 57.085 27.570 ;
        RECT 57.395 27.400 57.565 27.570 ;
        RECT 57.875 27.400 58.045 27.570 ;
        RECT 58.355 27.400 58.525 27.570 ;
        RECT 58.835 27.400 59.005 27.570 ;
        RECT 59.315 27.400 59.485 27.570 ;
        RECT 59.795 27.400 59.965 27.570 ;
        RECT 60.275 27.400 60.445 27.570 ;
        RECT 60.755 27.400 60.925 27.570 ;
        RECT 61.235 27.400 61.405 27.570 ;
        RECT 61.715 27.400 61.885 27.570 ;
        RECT 62.195 27.400 62.365 27.570 ;
        RECT 62.675 27.400 62.845 27.570 ;
        RECT 63.155 27.400 63.325 27.570 ;
        RECT 63.635 27.400 63.805 27.570 ;
        RECT 64.115 27.400 64.285 27.570 ;
        RECT 64.595 27.400 64.765 27.570 ;
        RECT 65.075 27.400 65.245 27.570 ;
        RECT 65.555 27.400 65.725 27.570 ;
        RECT 66.035 27.400 66.205 27.570 ;
        RECT 66.515 27.400 66.685 27.570 ;
        RECT 66.995 27.400 67.165 27.570 ;
        RECT 67.475 27.400 67.645 27.570 ;
        RECT 67.955 27.400 68.125 27.570 ;
        RECT 68.435 27.400 68.605 27.570 ;
        RECT 68.915 27.400 69.085 27.570 ;
        RECT 69.395 27.400 69.565 27.570 ;
        RECT 69.875 27.400 70.045 27.570 ;
        RECT 70.355 27.400 70.525 27.570 ;
        RECT 70.835 27.400 71.005 27.570 ;
        RECT 71.315 27.400 71.485 27.570 ;
        RECT 71.795 27.400 71.965 27.570 ;
        RECT 72.275 27.400 72.445 27.570 ;
        RECT 72.755 27.400 72.925 27.570 ;
      LAYER met1 ;
        RECT 0.000 37.210 88.240 38.650 ;
        RECT 0.000 26.865 88.240 28.305 ;
        RECT 0.000 3.220 88.240 11.220 ;
      LAYER via ;
        RECT 5.265 38.140 5.525 38.400 ;
        RECT 5.605 38.140 5.865 38.400 ;
        RECT 5.925 38.140 6.185 38.400 ;
        RECT 6.350 38.140 6.610 38.400 ;
        RECT 6.690 38.140 6.950 38.400 ;
        RECT 5.265 37.815 5.525 38.075 ;
        RECT 5.605 37.815 5.865 38.075 ;
        RECT 5.925 37.815 6.185 38.075 ;
        RECT 6.350 37.815 6.610 38.075 ;
        RECT 6.690 37.815 6.950 38.075 ;
        RECT 5.265 37.485 5.525 37.745 ;
        RECT 5.605 37.485 5.865 37.745 ;
        RECT 5.925 37.485 6.185 37.745 ;
        RECT 6.350 37.485 6.610 37.745 ;
        RECT 6.690 37.485 6.950 37.745 ;
        RECT 5.265 27.760 5.525 28.020 ;
        RECT 5.605 27.760 5.865 28.020 ;
        RECT 5.925 27.760 6.185 28.020 ;
        RECT 6.350 27.760 6.610 28.020 ;
        RECT 6.690 27.760 6.950 28.020 ;
        RECT 5.265 27.435 5.525 27.695 ;
        RECT 5.605 27.435 5.865 27.695 ;
        RECT 5.925 27.435 6.185 27.695 ;
        RECT 6.350 27.435 6.610 27.695 ;
        RECT 6.690 27.435 6.950 27.695 ;
        RECT 5.265 27.105 5.525 27.365 ;
        RECT 5.605 27.105 5.865 27.365 ;
        RECT 5.925 27.105 6.185 27.365 ;
        RECT 6.350 27.105 6.610 27.365 ;
        RECT 6.690 27.105 6.950 27.365 ;
        RECT 5.265 10.580 5.525 10.840 ;
        RECT 5.605 10.580 5.865 10.840 ;
        RECT 5.925 10.580 6.185 10.840 ;
        RECT 6.350 10.580 6.610 10.840 ;
        RECT 6.690 10.580 6.950 10.840 ;
        RECT 5.265 10.255 5.525 10.515 ;
        RECT 5.605 10.255 5.865 10.515 ;
        RECT 5.925 10.255 6.185 10.515 ;
        RECT 6.350 10.255 6.610 10.515 ;
        RECT 6.690 10.255 6.950 10.515 ;
        RECT 5.265 9.925 5.525 10.185 ;
        RECT 5.605 9.925 5.865 10.185 ;
        RECT 5.925 9.925 6.185 10.185 ;
        RECT 6.350 9.925 6.610 10.185 ;
        RECT 6.690 9.925 6.950 10.185 ;
        RECT 5.265 9.425 5.525 9.685 ;
        RECT 5.605 9.425 5.865 9.685 ;
        RECT 5.925 9.425 6.185 9.685 ;
        RECT 6.350 9.425 6.610 9.685 ;
        RECT 6.690 9.425 6.950 9.685 ;
        RECT 5.265 9.100 5.525 9.360 ;
        RECT 5.605 9.100 5.865 9.360 ;
        RECT 5.925 9.100 6.185 9.360 ;
        RECT 6.350 9.100 6.610 9.360 ;
        RECT 6.690 9.100 6.950 9.360 ;
        RECT 5.265 8.770 5.525 9.030 ;
        RECT 5.605 8.770 5.865 9.030 ;
        RECT 5.925 8.770 6.185 9.030 ;
        RECT 6.350 8.770 6.610 9.030 ;
        RECT 6.690 8.770 6.950 9.030 ;
        RECT 5.265 8.155 5.525 8.415 ;
        RECT 5.605 8.155 5.865 8.415 ;
        RECT 5.925 8.155 6.185 8.415 ;
        RECT 6.350 8.155 6.610 8.415 ;
        RECT 6.690 8.155 6.950 8.415 ;
        RECT 5.265 7.830 5.525 8.090 ;
        RECT 5.605 7.830 5.865 8.090 ;
        RECT 5.925 7.830 6.185 8.090 ;
        RECT 6.350 7.830 6.610 8.090 ;
        RECT 6.690 7.830 6.950 8.090 ;
        RECT 5.265 7.500 5.525 7.760 ;
        RECT 5.605 7.500 5.865 7.760 ;
        RECT 5.925 7.500 6.185 7.760 ;
        RECT 6.350 7.500 6.610 7.760 ;
        RECT 6.690 7.500 6.950 7.760 ;
        RECT 5.265 7.000 5.525 7.260 ;
        RECT 5.605 7.000 5.865 7.260 ;
        RECT 5.925 7.000 6.185 7.260 ;
        RECT 6.350 7.000 6.610 7.260 ;
        RECT 6.690 7.000 6.950 7.260 ;
        RECT 5.265 6.675 5.525 6.935 ;
        RECT 5.605 6.675 5.865 6.935 ;
        RECT 5.925 6.675 6.185 6.935 ;
        RECT 6.350 6.675 6.610 6.935 ;
        RECT 6.690 6.675 6.950 6.935 ;
        RECT 5.265 6.345 5.525 6.605 ;
        RECT 5.605 6.345 5.865 6.605 ;
        RECT 5.925 6.345 6.185 6.605 ;
        RECT 6.350 6.345 6.610 6.605 ;
        RECT 6.690 6.345 6.950 6.605 ;
        RECT 5.265 5.825 5.525 6.085 ;
        RECT 5.605 5.825 5.865 6.085 ;
        RECT 5.925 5.825 6.185 6.085 ;
        RECT 6.350 5.825 6.610 6.085 ;
        RECT 6.690 5.825 6.950 6.085 ;
        RECT 5.265 5.500 5.525 5.760 ;
        RECT 5.605 5.500 5.865 5.760 ;
        RECT 5.925 5.500 6.185 5.760 ;
        RECT 6.350 5.500 6.610 5.760 ;
        RECT 6.690 5.500 6.950 5.760 ;
        RECT 5.265 5.170 5.525 5.430 ;
        RECT 5.605 5.170 5.865 5.430 ;
        RECT 5.925 5.170 6.185 5.430 ;
        RECT 6.350 5.170 6.610 5.430 ;
        RECT 6.690 5.170 6.950 5.430 ;
        RECT 5.265 4.670 5.525 4.930 ;
        RECT 5.605 4.670 5.865 4.930 ;
        RECT 5.925 4.670 6.185 4.930 ;
        RECT 6.350 4.670 6.610 4.930 ;
        RECT 6.690 4.670 6.950 4.930 ;
        RECT 5.265 4.345 5.525 4.605 ;
        RECT 5.605 4.345 5.865 4.605 ;
        RECT 5.925 4.345 6.185 4.605 ;
        RECT 6.350 4.345 6.610 4.605 ;
        RECT 6.690 4.345 6.950 4.605 ;
        RECT 5.265 4.015 5.525 4.275 ;
        RECT 5.605 4.015 5.865 4.275 ;
        RECT 5.925 4.015 6.185 4.275 ;
        RECT 6.350 4.015 6.610 4.275 ;
        RECT 6.690 4.015 6.950 4.275 ;
      LAYER met2 ;
        RECT 5.085 3.600 7.085 38.865 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 7.740 46.230 81.240 47.660 ;
        RECT 7.740 18.355 9.170 46.230 ;
        RECT 14.675 39.715 63.815 41.320 ;
        RECT 54.990 30.975 73.410 31.970 ;
        RECT 12.600 29.370 73.410 30.975 ;
        RECT 79.810 18.355 81.240 46.230 ;
        RECT 7.740 16.925 81.240 18.355 ;
      LAYER li1 ;
        RECT 8.425 41.045 80.555 46.975 ;
        RECT 8.425 21.745 12.455 41.045 ;
        RECT 14.950 39.880 15.240 41.045 ;
        RECT 15.680 40.245 15.930 41.045 ;
        RECT 16.600 40.245 16.770 41.045 ;
        RECT 17.440 40.245 17.610 41.045 ;
        RECT 18.280 40.245 18.450 41.045 ;
        RECT 19.120 39.905 19.375 41.045 ;
        RECT 21.435 39.905 21.700 41.045 ;
        RECT 22.370 40.245 22.540 41.045 ;
        RECT 23.210 40.585 23.420 41.045 ;
        RECT 25.530 39.880 25.820 41.045 ;
        RECT 27.930 40.585 28.140 41.045 ;
        RECT 28.810 40.245 28.980 41.045 ;
        RECT 29.650 39.905 29.915 41.045 ;
        RECT 31.975 39.905 32.230 41.045 ;
        RECT 32.900 40.245 33.070 41.045 ;
        RECT 33.740 40.245 33.910 41.045 ;
        RECT 34.580 40.245 34.750 41.045 ;
        RECT 35.420 40.245 35.670 41.045 ;
        RECT 36.210 40.585 36.420 41.045 ;
        RECT 37.090 40.245 37.260 41.045 ;
        RECT 37.930 39.905 38.195 41.045 ;
        RECT 40.520 40.245 40.770 41.045 ;
        RECT 41.440 40.245 41.610 41.045 ;
        RECT 42.280 40.245 42.450 41.045 ;
        RECT 43.120 40.245 43.290 41.045 ;
        RECT 43.960 39.905 44.215 41.045 ;
        RECT 44.390 39.880 44.680 41.045 ;
        RECT 46.790 40.585 47.000 41.045 ;
        RECT 47.670 40.245 47.840 41.045 ;
        RECT 48.510 39.905 48.775 41.045 ;
        RECT 50.835 39.905 51.090 41.045 ;
        RECT 51.760 40.245 51.930 41.045 ;
        RECT 52.600 40.245 52.770 41.045 ;
        RECT 53.440 40.245 53.610 41.045 ;
        RECT 54.280 40.245 54.530 41.045 ;
        RECT 55.070 40.585 55.280 41.045 ;
        RECT 55.950 40.245 56.120 41.045 ;
        RECT 56.790 39.905 57.055 41.045 ;
        RECT 59.115 39.905 59.370 41.045 ;
        RECT 60.040 40.245 60.210 41.045 ;
        RECT 60.880 40.245 61.050 41.045 ;
        RECT 61.720 40.245 61.890 41.045 ;
        RECT 62.560 40.245 62.810 41.045 ;
        RECT 63.250 39.880 63.540 41.045 ;
        RECT 55.320 31.470 73.080 31.640 ;
        RECT 12.790 30.700 54.650 30.870 ;
        RECT 12.875 29.535 13.165 30.700 ;
        RECT 15.275 30.240 15.485 30.700 ;
        RECT 16.155 29.900 16.325 30.700 ;
        RECT 16.995 29.560 17.260 30.700 ;
        RECT 21.745 29.900 21.995 30.700 ;
        RECT 22.505 29.900 22.835 30.700 ;
        RECT 25.395 30.240 25.605 30.700 ;
        RECT 26.275 29.900 26.445 30.700 ;
        RECT 27.115 29.560 27.380 30.700 ;
        RECT 29.435 29.535 29.725 30.700 ;
        RECT 31.835 30.240 32.045 30.700 ;
        RECT 32.715 29.900 32.885 30.700 ;
        RECT 33.555 29.560 33.820 30.700 ;
        RECT 38.305 29.900 38.555 30.700 ;
        RECT 39.065 29.900 39.395 30.700 ;
        RECT 40.015 29.535 40.305 30.700 ;
        RECT 46.095 30.240 46.305 30.700 ;
        RECT 46.975 29.900 47.145 30.700 ;
        RECT 47.815 29.560 48.080 30.700 ;
        RECT 52.565 29.900 52.815 30.700 ;
        RECT 53.325 29.900 53.655 30.700 ;
        RECT 54.275 29.535 54.565 30.700 ;
        RECT 55.480 29.660 56.010 31.240 ;
        RECT 56.760 29.660 57.650 31.240 ;
        RECT 58.320 29.660 59.210 31.240 ;
        RECT 59.880 29.660 60.770 31.240 ;
        RECT 61.440 29.660 62.330 31.240 ;
        RECT 63.000 29.660 63.890 31.240 ;
        RECT 64.560 29.660 65.450 31.240 ;
        RECT 66.120 29.660 67.010 31.240 ;
        RECT 67.730 29.930 68.620 31.160 ;
        RECT 69.310 29.930 70.200 31.160 ;
        RECT 70.850 29.930 71.740 31.160 ;
        RECT 72.400 29.660 72.970 31.240 ;
        RECT 75.225 21.745 80.555 41.045 ;
        RECT 8.425 17.610 80.555 21.745 ;
      LAYER mcon ;
        RECT 9.205 41.695 9.375 41.865 ;
        RECT 9.565 41.695 9.735 41.865 ;
        RECT 9.925 41.695 10.095 41.865 ;
        RECT 10.285 41.695 10.455 41.865 ;
        RECT 10.645 41.695 10.815 41.865 ;
        RECT 11.005 41.695 11.175 41.865 ;
        RECT 11.365 41.695 11.535 41.865 ;
        RECT 11.725 41.695 11.895 41.865 ;
        RECT 12.085 41.695 12.255 41.865 ;
        RECT 76.360 41.695 76.530 41.865 ;
        RECT 76.720 41.695 76.890 41.865 ;
        RECT 77.080 41.695 77.250 41.865 ;
        RECT 77.440 41.695 77.610 41.865 ;
        RECT 77.800 41.695 77.970 41.865 ;
        RECT 78.160 41.695 78.330 41.865 ;
        RECT 78.520 41.695 78.690 41.865 ;
        RECT 78.880 41.695 79.050 41.865 ;
        RECT 79.240 41.695 79.410 41.865 ;
        RECT 9.205 41.180 9.375 41.350 ;
        RECT 9.565 41.180 9.735 41.350 ;
        RECT 9.925 41.180 10.095 41.350 ;
        RECT 10.285 41.180 10.455 41.350 ;
        RECT 10.645 41.180 10.815 41.350 ;
        RECT 11.005 41.180 11.175 41.350 ;
        RECT 11.365 41.180 11.535 41.350 ;
        RECT 11.725 41.180 11.895 41.350 ;
        RECT 12.085 41.180 12.255 41.350 ;
        RECT 15.010 41.045 15.180 41.215 ;
        RECT 15.470 41.045 15.640 41.215 ;
        RECT 15.930 41.045 16.100 41.215 ;
        RECT 16.390 41.045 16.560 41.215 ;
        RECT 16.850 41.045 17.020 41.215 ;
        RECT 17.310 41.045 17.480 41.215 ;
        RECT 17.770 41.045 17.940 41.215 ;
        RECT 18.230 41.045 18.400 41.215 ;
        RECT 18.690 41.045 18.860 41.215 ;
        RECT 19.150 41.045 19.320 41.215 ;
        RECT 19.610 41.045 19.780 41.215 ;
        RECT 20.070 41.045 20.240 41.215 ;
        RECT 20.530 41.045 20.700 41.215 ;
        RECT 20.990 41.045 21.160 41.215 ;
        RECT 21.450 41.045 21.620 41.215 ;
        RECT 21.910 41.045 22.080 41.215 ;
        RECT 22.370 41.045 22.540 41.215 ;
        RECT 22.830 41.045 23.000 41.215 ;
        RECT 23.290 41.045 23.460 41.215 ;
        RECT 23.750 41.045 23.920 41.215 ;
        RECT 24.210 41.045 24.380 41.215 ;
        RECT 24.670 41.045 24.840 41.215 ;
        RECT 25.130 41.045 25.300 41.215 ;
        RECT 25.590 41.045 25.760 41.215 ;
        RECT 26.050 41.045 26.220 41.215 ;
        RECT 26.510 41.045 26.680 41.215 ;
        RECT 26.970 41.045 27.140 41.215 ;
        RECT 27.430 41.045 27.600 41.215 ;
        RECT 27.890 41.045 28.060 41.215 ;
        RECT 28.350 41.045 28.520 41.215 ;
        RECT 28.810 41.045 28.980 41.215 ;
        RECT 29.270 41.045 29.440 41.215 ;
        RECT 29.730 41.045 29.900 41.215 ;
        RECT 30.190 41.045 30.360 41.215 ;
        RECT 30.650 41.045 30.820 41.215 ;
        RECT 31.110 41.045 31.280 41.215 ;
        RECT 31.570 41.045 31.740 41.215 ;
        RECT 32.030 41.045 32.200 41.215 ;
        RECT 32.490 41.045 32.660 41.215 ;
        RECT 32.950 41.045 33.120 41.215 ;
        RECT 33.410 41.045 33.580 41.215 ;
        RECT 33.870 41.045 34.040 41.215 ;
        RECT 34.330 41.045 34.500 41.215 ;
        RECT 34.790 41.045 34.960 41.215 ;
        RECT 35.250 41.045 35.420 41.215 ;
        RECT 35.710 41.045 35.880 41.215 ;
        RECT 36.170 41.045 36.340 41.215 ;
        RECT 36.630 41.045 36.800 41.215 ;
        RECT 37.090 41.045 37.260 41.215 ;
        RECT 37.550 41.045 37.720 41.215 ;
        RECT 38.010 41.045 38.180 41.215 ;
        RECT 38.470 41.045 38.640 41.215 ;
        RECT 38.930 41.045 39.100 41.215 ;
        RECT 39.390 41.045 39.560 41.215 ;
        RECT 39.850 41.045 40.020 41.215 ;
        RECT 40.310 41.045 40.480 41.215 ;
        RECT 40.770 41.045 40.940 41.215 ;
        RECT 41.230 41.045 41.400 41.215 ;
        RECT 41.690 41.045 41.860 41.215 ;
        RECT 42.150 41.045 42.320 41.215 ;
        RECT 42.610 41.045 42.780 41.215 ;
        RECT 43.070 41.045 43.240 41.215 ;
        RECT 43.530 41.045 43.700 41.215 ;
        RECT 43.990 41.045 44.160 41.215 ;
        RECT 44.450 41.045 44.620 41.215 ;
        RECT 44.910 41.045 45.080 41.215 ;
        RECT 45.370 41.045 45.540 41.215 ;
        RECT 45.830 41.045 46.000 41.215 ;
        RECT 46.290 41.045 46.460 41.215 ;
        RECT 46.750 41.045 46.920 41.215 ;
        RECT 47.210 41.045 47.380 41.215 ;
        RECT 47.670 41.045 47.840 41.215 ;
        RECT 48.130 41.045 48.300 41.215 ;
        RECT 48.590 41.045 48.760 41.215 ;
        RECT 49.050 41.045 49.220 41.215 ;
        RECT 49.510 41.045 49.680 41.215 ;
        RECT 49.970 41.045 50.140 41.215 ;
        RECT 50.430 41.045 50.600 41.215 ;
        RECT 50.890 41.045 51.060 41.215 ;
        RECT 51.350 41.045 51.520 41.215 ;
        RECT 51.810 41.045 51.980 41.215 ;
        RECT 52.270 41.045 52.440 41.215 ;
        RECT 52.730 41.045 52.900 41.215 ;
        RECT 53.190 41.045 53.360 41.215 ;
        RECT 53.650 41.045 53.820 41.215 ;
        RECT 54.110 41.045 54.280 41.215 ;
        RECT 54.570 41.045 54.740 41.215 ;
        RECT 55.030 41.045 55.200 41.215 ;
        RECT 55.490 41.045 55.660 41.215 ;
        RECT 55.950 41.045 56.120 41.215 ;
        RECT 56.410 41.045 56.580 41.215 ;
        RECT 56.870 41.045 57.040 41.215 ;
        RECT 57.330 41.045 57.500 41.215 ;
        RECT 57.790 41.045 57.960 41.215 ;
        RECT 58.250 41.045 58.420 41.215 ;
        RECT 58.710 41.045 58.880 41.215 ;
        RECT 59.170 41.045 59.340 41.215 ;
        RECT 59.630 41.045 59.800 41.215 ;
        RECT 60.090 41.045 60.260 41.215 ;
        RECT 60.550 41.045 60.720 41.215 ;
        RECT 61.010 41.045 61.180 41.215 ;
        RECT 61.470 41.045 61.640 41.215 ;
        RECT 61.930 41.045 62.100 41.215 ;
        RECT 62.390 41.045 62.560 41.215 ;
        RECT 62.850 41.045 63.020 41.215 ;
        RECT 63.310 41.045 63.480 41.215 ;
        RECT 76.360 41.180 76.530 41.350 ;
        RECT 76.720 41.180 76.890 41.350 ;
        RECT 77.080 41.180 77.250 41.350 ;
        RECT 77.440 41.180 77.610 41.350 ;
        RECT 77.800 41.180 77.970 41.350 ;
        RECT 78.160 41.180 78.330 41.350 ;
        RECT 78.520 41.180 78.690 41.350 ;
        RECT 78.880 41.180 79.050 41.350 ;
        RECT 79.240 41.180 79.410 41.350 ;
        RECT 9.175 31.465 9.345 31.635 ;
        RECT 9.535 31.465 9.705 31.635 ;
        RECT 9.895 31.465 10.065 31.635 ;
        RECT 10.255 31.465 10.425 31.635 ;
        RECT 10.615 31.465 10.785 31.635 ;
        RECT 10.975 31.465 11.145 31.635 ;
        RECT 11.335 31.465 11.505 31.635 ;
        RECT 11.695 31.465 11.865 31.635 ;
        RECT 12.055 31.465 12.225 31.635 ;
        RECT 55.475 31.470 55.645 31.640 ;
        RECT 55.955 31.470 56.125 31.640 ;
        RECT 56.435 31.470 56.605 31.640 ;
        RECT 56.915 31.470 57.085 31.640 ;
        RECT 57.395 31.470 57.565 31.640 ;
        RECT 57.875 31.470 58.045 31.640 ;
        RECT 58.355 31.470 58.525 31.640 ;
        RECT 58.835 31.470 59.005 31.640 ;
        RECT 59.315 31.470 59.485 31.640 ;
        RECT 59.795 31.470 59.965 31.640 ;
        RECT 60.275 31.470 60.445 31.640 ;
        RECT 60.755 31.470 60.925 31.640 ;
        RECT 61.235 31.470 61.405 31.640 ;
        RECT 61.715 31.470 61.885 31.640 ;
        RECT 62.195 31.470 62.365 31.640 ;
        RECT 62.675 31.470 62.845 31.640 ;
        RECT 63.155 31.470 63.325 31.640 ;
        RECT 63.635 31.470 63.805 31.640 ;
        RECT 64.115 31.470 64.285 31.640 ;
        RECT 64.595 31.470 64.765 31.640 ;
        RECT 65.075 31.470 65.245 31.640 ;
        RECT 65.555 31.470 65.725 31.640 ;
        RECT 66.035 31.470 66.205 31.640 ;
        RECT 66.515 31.470 66.685 31.640 ;
        RECT 66.995 31.470 67.165 31.640 ;
        RECT 67.475 31.470 67.645 31.640 ;
        RECT 67.955 31.470 68.125 31.640 ;
        RECT 68.435 31.470 68.605 31.640 ;
        RECT 68.915 31.470 69.085 31.640 ;
        RECT 69.395 31.470 69.565 31.640 ;
        RECT 69.875 31.470 70.045 31.640 ;
        RECT 70.355 31.470 70.525 31.640 ;
        RECT 70.835 31.470 71.005 31.640 ;
        RECT 71.315 31.470 71.485 31.640 ;
        RECT 71.795 31.470 71.965 31.640 ;
        RECT 72.275 31.470 72.445 31.640 ;
        RECT 72.755 31.470 72.925 31.640 ;
        RECT 76.330 31.465 76.500 31.635 ;
        RECT 76.690 31.465 76.860 31.635 ;
        RECT 77.050 31.465 77.220 31.635 ;
        RECT 77.410 31.465 77.580 31.635 ;
        RECT 77.770 31.465 77.940 31.635 ;
        RECT 78.130 31.465 78.300 31.635 ;
        RECT 78.490 31.465 78.660 31.635 ;
        RECT 78.850 31.465 79.020 31.635 ;
        RECT 79.210 31.465 79.380 31.635 ;
        RECT 9.175 30.950 9.345 31.120 ;
        RECT 9.535 30.950 9.705 31.120 ;
        RECT 9.895 30.950 10.065 31.120 ;
        RECT 10.255 30.950 10.425 31.120 ;
        RECT 10.615 30.950 10.785 31.120 ;
        RECT 10.975 30.950 11.145 31.120 ;
        RECT 11.335 30.950 11.505 31.120 ;
        RECT 11.695 30.950 11.865 31.120 ;
        RECT 12.055 30.950 12.225 31.120 ;
        RECT 55.480 30.960 55.650 31.130 ;
        RECT 55.840 30.960 56.010 31.130 ;
        RECT 12.935 30.700 13.105 30.870 ;
        RECT 13.395 30.700 13.565 30.870 ;
        RECT 13.855 30.700 14.025 30.870 ;
        RECT 14.315 30.700 14.485 30.870 ;
        RECT 14.775 30.700 14.945 30.870 ;
        RECT 15.235 30.700 15.405 30.870 ;
        RECT 15.695 30.700 15.865 30.870 ;
        RECT 16.155 30.700 16.325 30.870 ;
        RECT 16.615 30.700 16.785 30.870 ;
        RECT 17.075 30.700 17.245 30.870 ;
        RECT 17.535 30.700 17.705 30.870 ;
        RECT 17.995 30.700 18.165 30.870 ;
        RECT 18.455 30.700 18.625 30.870 ;
        RECT 18.915 30.700 19.085 30.870 ;
        RECT 19.375 30.700 19.545 30.870 ;
        RECT 19.835 30.700 20.005 30.870 ;
        RECT 20.295 30.700 20.465 30.870 ;
        RECT 20.755 30.700 20.925 30.870 ;
        RECT 21.215 30.700 21.385 30.870 ;
        RECT 21.675 30.700 21.845 30.870 ;
        RECT 22.135 30.700 22.305 30.870 ;
        RECT 22.595 30.700 22.765 30.870 ;
        RECT 23.055 30.700 23.225 30.870 ;
        RECT 23.515 30.700 23.685 30.870 ;
        RECT 23.975 30.700 24.145 30.870 ;
        RECT 24.435 30.700 24.605 30.870 ;
        RECT 24.895 30.700 25.065 30.870 ;
        RECT 25.355 30.700 25.525 30.870 ;
        RECT 25.815 30.700 25.985 30.870 ;
        RECT 26.275 30.700 26.445 30.870 ;
        RECT 26.735 30.700 26.905 30.870 ;
        RECT 27.195 30.700 27.365 30.870 ;
        RECT 27.655 30.700 27.825 30.870 ;
        RECT 28.115 30.700 28.285 30.870 ;
        RECT 28.575 30.700 28.745 30.870 ;
        RECT 29.035 30.700 29.205 30.870 ;
        RECT 29.495 30.700 29.665 30.870 ;
        RECT 29.955 30.700 30.125 30.870 ;
        RECT 30.415 30.700 30.585 30.870 ;
        RECT 30.875 30.700 31.045 30.870 ;
        RECT 31.335 30.700 31.505 30.870 ;
        RECT 31.795 30.700 31.965 30.870 ;
        RECT 32.255 30.700 32.425 30.870 ;
        RECT 32.715 30.700 32.885 30.870 ;
        RECT 33.175 30.700 33.345 30.870 ;
        RECT 33.635 30.700 33.805 30.870 ;
        RECT 34.095 30.700 34.265 30.870 ;
        RECT 34.555 30.700 34.725 30.870 ;
        RECT 35.015 30.700 35.185 30.870 ;
        RECT 35.475 30.700 35.645 30.870 ;
        RECT 35.935 30.700 36.105 30.870 ;
        RECT 36.395 30.700 36.565 30.870 ;
        RECT 36.855 30.700 37.025 30.870 ;
        RECT 37.315 30.700 37.485 30.870 ;
        RECT 37.775 30.700 37.945 30.870 ;
        RECT 38.235 30.700 38.405 30.870 ;
        RECT 38.695 30.700 38.865 30.870 ;
        RECT 39.155 30.700 39.325 30.870 ;
        RECT 39.615 30.700 39.785 30.870 ;
        RECT 40.075 30.700 40.245 30.870 ;
        RECT 40.535 30.700 40.705 30.870 ;
        RECT 40.995 30.700 41.165 30.870 ;
        RECT 41.455 30.700 41.625 30.870 ;
        RECT 41.915 30.700 42.085 30.870 ;
        RECT 42.375 30.700 42.545 30.870 ;
        RECT 42.835 30.700 43.005 30.870 ;
        RECT 43.295 30.700 43.465 30.870 ;
        RECT 43.755 30.700 43.925 30.870 ;
        RECT 44.215 30.700 44.385 30.870 ;
        RECT 44.675 30.700 44.845 30.870 ;
        RECT 45.135 30.700 45.305 30.870 ;
        RECT 45.595 30.700 45.765 30.870 ;
        RECT 46.055 30.700 46.225 30.870 ;
        RECT 46.515 30.700 46.685 30.870 ;
        RECT 46.975 30.700 47.145 30.870 ;
        RECT 47.435 30.700 47.605 30.870 ;
        RECT 47.895 30.700 48.065 30.870 ;
        RECT 48.355 30.700 48.525 30.870 ;
        RECT 48.815 30.700 48.985 30.870 ;
        RECT 49.275 30.700 49.445 30.870 ;
        RECT 49.735 30.700 49.905 30.870 ;
        RECT 50.195 30.700 50.365 30.870 ;
        RECT 50.655 30.700 50.825 30.870 ;
        RECT 51.115 30.700 51.285 30.870 ;
        RECT 51.575 30.700 51.745 30.870 ;
        RECT 52.035 30.700 52.205 30.870 ;
        RECT 52.495 30.700 52.665 30.870 ;
        RECT 52.955 30.700 53.125 30.870 ;
        RECT 53.415 30.700 53.585 30.870 ;
        RECT 53.875 30.700 54.045 30.870 ;
        RECT 54.335 30.700 54.505 30.870 ;
        RECT 56.760 30.960 56.930 31.130 ;
        RECT 57.120 30.960 57.290 31.130 ;
        RECT 57.480 30.960 57.650 31.130 ;
        RECT 58.320 30.960 58.490 31.130 ;
        RECT 58.680 30.960 58.850 31.130 ;
        RECT 59.040 30.960 59.210 31.130 ;
        RECT 59.880 30.960 60.050 31.130 ;
        RECT 60.240 30.960 60.410 31.130 ;
        RECT 60.600 30.960 60.770 31.130 ;
        RECT 61.440 30.960 61.610 31.130 ;
        RECT 61.800 30.960 61.970 31.130 ;
        RECT 62.160 30.960 62.330 31.130 ;
        RECT 63.000 30.960 63.170 31.130 ;
        RECT 63.360 30.960 63.530 31.130 ;
        RECT 63.720 30.960 63.890 31.130 ;
        RECT 64.560 30.960 64.730 31.130 ;
        RECT 64.920 30.960 65.090 31.130 ;
        RECT 65.280 30.960 65.450 31.130 ;
        RECT 66.120 30.960 66.290 31.130 ;
        RECT 66.480 30.960 66.650 31.130 ;
        RECT 66.840 30.960 67.010 31.130 ;
        RECT 67.730 30.960 67.900 31.130 ;
        RECT 68.090 30.960 68.260 31.130 ;
        RECT 68.450 30.960 68.620 31.130 ;
        RECT 69.310 30.960 69.480 31.130 ;
        RECT 69.670 30.960 69.840 31.130 ;
        RECT 70.030 30.960 70.200 31.130 ;
        RECT 70.850 30.960 71.020 31.130 ;
        RECT 71.210 30.960 71.380 31.130 ;
        RECT 71.570 30.960 71.740 31.130 ;
        RECT 72.400 30.960 72.570 31.130 ;
        RECT 72.760 30.960 72.930 31.130 ;
        RECT 76.330 30.950 76.500 31.120 ;
        RECT 76.690 30.950 76.860 31.120 ;
        RECT 77.050 30.950 77.220 31.120 ;
        RECT 77.410 30.950 77.580 31.120 ;
        RECT 77.770 30.950 77.940 31.120 ;
        RECT 78.130 30.950 78.300 31.120 ;
        RECT 78.490 30.950 78.660 31.120 ;
        RECT 78.850 30.950 79.020 31.120 ;
        RECT 79.210 30.950 79.380 31.120 ;
        RECT 10.585 20.065 10.755 20.235 ;
        RECT 10.945 20.065 11.115 20.235 ;
        RECT 11.305 20.065 11.475 20.235 ;
        RECT 11.665 20.065 11.835 20.235 ;
        RECT 12.025 20.065 12.195 20.235 ;
        RECT 12.385 20.065 12.555 20.235 ;
        RECT 12.745 20.065 12.915 20.235 ;
        RECT 13.105 20.065 13.275 20.235 ;
        RECT 13.465 20.065 13.635 20.235 ;
        RECT 14.150 20.065 14.320 20.235 ;
        RECT 14.510 20.065 14.680 20.235 ;
        RECT 14.870 20.065 15.040 20.235 ;
        RECT 15.230 20.065 15.400 20.235 ;
        RECT 15.590 20.065 15.760 20.235 ;
        RECT 15.950 20.065 16.120 20.235 ;
        RECT 16.310 20.065 16.480 20.235 ;
        RECT 16.670 20.065 16.840 20.235 ;
        RECT 17.030 20.065 17.200 20.235 ;
        RECT 17.835 20.065 18.005 20.235 ;
        RECT 18.195 20.065 18.365 20.235 ;
        RECT 18.555 20.065 18.725 20.235 ;
        RECT 18.915 20.065 19.085 20.235 ;
        RECT 19.275 20.065 19.445 20.235 ;
        RECT 19.635 20.065 19.805 20.235 ;
        RECT 19.995 20.065 20.165 20.235 ;
        RECT 20.355 20.065 20.525 20.235 ;
        RECT 20.715 20.065 20.885 20.235 ;
        RECT 21.400 20.065 21.570 20.235 ;
        RECT 21.760 20.065 21.930 20.235 ;
        RECT 22.120 20.065 22.290 20.235 ;
        RECT 22.480 20.065 22.650 20.235 ;
        RECT 22.840 20.065 23.010 20.235 ;
        RECT 23.200 20.065 23.370 20.235 ;
        RECT 23.560 20.065 23.730 20.235 ;
        RECT 23.920 20.065 24.090 20.235 ;
        RECT 24.280 20.065 24.450 20.235 ;
        RECT 25.460 20.065 25.630 20.235 ;
        RECT 25.820 20.065 25.990 20.235 ;
        RECT 26.180 20.065 26.350 20.235 ;
        RECT 26.540 20.065 26.710 20.235 ;
        RECT 26.900 20.065 27.070 20.235 ;
        RECT 27.260 20.065 27.430 20.235 ;
        RECT 27.620 20.065 27.790 20.235 ;
        RECT 27.980 20.065 28.150 20.235 ;
        RECT 28.340 20.065 28.510 20.235 ;
        RECT 29.025 20.065 29.195 20.235 ;
        RECT 29.385 20.065 29.555 20.235 ;
        RECT 29.745 20.065 29.915 20.235 ;
        RECT 30.105 20.065 30.275 20.235 ;
        RECT 30.465 20.065 30.635 20.235 ;
        RECT 30.825 20.065 30.995 20.235 ;
        RECT 31.185 20.065 31.355 20.235 ;
        RECT 31.545 20.065 31.715 20.235 ;
        RECT 31.905 20.065 32.075 20.235 ;
        RECT 32.710 20.065 32.880 20.235 ;
        RECT 33.070 20.065 33.240 20.235 ;
        RECT 33.430 20.065 33.600 20.235 ;
        RECT 33.790 20.065 33.960 20.235 ;
        RECT 34.150 20.065 34.320 20.235 ;
        RECT 34.510 20.065 34.680 20.235 ;
        RECT 34.870 20.065 35.040 20.235 ;
        RECT 35.230 20.065 35.400 20.235 ;
        RECT 35.590 20.065 35.760 20.235 ;
        RECT 36.275 20.065 36.445 20.235 ;
        RECT 36.635 20.065 36.805 20.235 ;
        RECT 36.995 20.065 37.165 20.235 ;
        RECT 37.355 20.065 37.525 20.235 ;
        RECT 37.715 20.065 37.885 20.235 ;
        RECT 38.075 20.065 38.245 20.235 ;
        RECT 38.435 20.065 38.605 20.235 ;
        RECT 38.795 20.065 38.965 20.235 ;
        RECT 39.155 20.065 39.325 20.235 ;
        RECT 40.390 20.065 40.560 20.235 ;
        RECT 40.750 20.065 40.920 20.235 ;
        RECT 41.110 20.065 41.280 20.235 ;
        RECT 41.470 20.065 41.640 20.235 ;
        RECT 41.830 20.065 42.000 20.235 ;
        RECT 42.190 20.065 42.360 20.235 ;
        RECT 42.550 20.065 42.720 20.235 ;
        RECT 42.910 20.065 43.080 20.235 ;
        RECT 43.270 20.065 43.440 20.235 ;
        RECT 43.955 20.065 44.125 20.235 ;
        RECT 44.315 20.065 44.485 20.235 ;
        RECT 44.675 20.065 44.845 20.235 ;
        RECT 45.035 20.065 45.205 20.235 ;
        RECT 45.395 20.065 45.565 20.235 ;
        RECT 45.755 20.065 45.925 20.235 ;
        RECT 46.115 20.065 46.285 20.235 ;
        RECT 46.475 20.065 46.645 20.235 ;
        RECT 46.835 20.065 47.005 20.235 ;
        RECT 47.640 20.065 47.810 20.235 ;
        RECT 48.000 20.065 48.170 20.235 ;
        RECT 48.360 20.065 48.530 20.235 ;
        RECT 48.720 20.065 48.890 20.235 ;
        RECT 49.080 20.065 49.250 20.235 ;
        RECT 49.440 20.065 49.610 20.235 ;
        RECT 49.800 20.065 49.970 20.235 ;
        RECT 50.160 20.065 50.330 20.235 ;
        RECT 50.520 20.065 50.690 20.235 ;
        RECT 51.205 20.065 51.375 20.235 ;
        RECT 51.565 20.065 51.735 20.235 ;
        RECT 51.925 20.065 52.095 20.235 ;
        RECT 52.285 20.065 52.455 20.235 ;
        RECT 52.645 20.065 52.815 20.235 ;
        RECT 53.005 20.065 53.175 20.235 ;
        RECT 53.365 20.065 53.535 20.235 ;
        RECT 53.725 20.065 53.895 20.235 ;
        RECT 54.085 20.065 54.255 20.235 ;
        RECT 55.265 20.065 55.435 20.235 ;
        RECT 55.625 20.065 55.795 20.235 ;
        RECT 55.985 20.065 56.155 20.235 ;
        RECT 56.345 20.065 56.515 20.235 ;
        RECT 56.705 20.065 56.875 20.235 ;
        RECT 57.065 20.065 57.235 20.235 ;
        RECT 57.425 20.065 57.595 20.235 ;
        RECT 57.785 20.065 57.955 20.235 ;
        RECT 58.145 20.065 58.315 20.235 ;
        RECT 58.830 20.065 59.000 20.235 ;
        RECT 59.190 20.065 59.360 20.235 ;
        RECT 59.550 20.065 59.720 20.235 ;
        RECT 59.910 20.065 60.080 20.235 ;
        RECT 60.270 20.065 60.440 20.235 ;
        RECT 60.630 20.065 60.800 20.235 ;
        RECT 60.990 20.065 61.160 20.235 ;
        RECT 61.350 20.065 61.520 20.235 ;
        RECT 61.710 20.065 61.880 20.235 ;
        RECT 62.515 20.065 62.685 20.235 ;
        RECT 62.875 20.065 63.045 20.235 ;
        RECT 63.235 20.065 63.405 20.235 ;
        RECT 63.595 20.065 63.765 20.235 ;
        RECT 63.955 20.065 64.125 20.235 ;
        RECT 64.315 20.065 64.485 20.235 ;
        RECT 64.675 20.065 64.845 20.235 ;
        RECT 65.035 20.065 65.205 20.235 ;
        RECT 65.395 20.065 65.565 20.235 ;
        RECT 66.080 20.065 66.250 20.235 ;
        RECT 66.440 20.065 66.610 20.235 ;
        RECT 66.800 20.065 66.970 20.235 ;
        RECT 67.160 20.065 67.330 20.235 ;
        RECT 67.520 20.065 67.690 20.235 ;
        RECT 67.880 20.065 68.050 20.235 ;
        RECT 68.240 20.065 68.410 20.235 ;
        RECT 68.600 20.065 68.770 20.235 ;
        RECT 68.960 20.065 69.130 20.235 ;
        RECT 70.010 20.065 70.180 20.235 ;
        RECT 70.370 20.065 70.540 20.235 ;
        RECT 70.730 20.065 70.900 20.235 ;
        RECT 71.090 20.065 71.260 20.235 ;
        RECT 71.450 20.065 71.620 20.235 ;
        RECT 71.810 20.065 71.980 20.235 ;
        RECT 72.170 20.065 72.340 20.235 ;
        RECT 72.530 20.065 72.700 20.235 ;
        RECT 72.890 20.065 73.060 20.235 ;
        RECT 73.575 20.065 73.745 20.235 ;
        RECT 73.935 20.065 74.105 20.235 ;
        RECT 74.295 20.065 74.465 20.235 ;
        RECT 74.655 20.065 74.825 20.235 ;
        RECT 75.015 20.065 75.185 20.235 ;
        RECT 75.375 20.065 75.545 20.235 ;
        RECT 75.735 20.065 75.905 20.235 ;
        RECT 76.095 20.065 76.265 20.235 ;
        RECT 76.455 20.065 76.625 20.235 ;
        RECT 10.585 19.550 10.755 19.720 ;
        RECT 10.945 19.550 11.115 19.720 ;
        RECT 11.305 19.550 11.475 19.720 ;
        RECT 11.665 19.550 11.835 19.720 ;
        RECT 12.025 19.550 12.195 19.720 ;
        RECT 12.385 19.550 12.555 19.720 ;
        RECT 12.745 19.550 12.915 19.720 ;
        RECT 13.105 19.550 13.275 19.720 ;
        RECT 13.465 19.550 13.635 19.720 ;
        RECT 14.150 19.550 14.320 19.720 ;
        RECT 14.510 19.550 14.680 19.720 ;
        RECT 14.870 19.550 15.040 19.720 ;
        RECT 15.230 19.550 15.400 19.720 ;
        RECT 15.590 19.550 15.760 19.720 ;
        RECT 15.950 19.550 16.120 19.720 ;
        RECT 16.310 19.550 16.480 19.720 ;
        RECT 16.670 19.550 16.840 19.720 ;
        RECT 17.030 19.550 17.200 19.720 ;
        RECT 17.835 19.550 18.005 19.720 ;
        RECT 18.195 19.550 18.365 19.720 ;
        RECT 18.555 19.550 18.725 19.720 ;
        RECT 18.915 19.550 19.085 19.720 ;
        RECT 19.275 19.550 19.445 19.720 ;
        RECT 19.635 19.550 19.805 19.720 ;
        RECT 19.995 19.550 20.165 19.720 ;
        RECT 20.355 19.550 20.525 19.720 ;
        RECT 20.715 19.550 20.885 19.720 ;
        RECT 21.400 19.550 21.570 19.720 ;
        RECT 21.760 19.550 21.930 19.720 ;
        RECT 22.120 19.550 22.290 19.720 ;
        RECT 22.480 19.550 22.650 19.720 ;
        RECT 22.840 19.550 23.010 19.720 ;
        RECT 23.200 19.550 23.370 19.720 ;
        RECT 23.560 19.550 23.730 19.720 ;
        RECT 23.920 19.550 24.090 19.720 ;
        RECT 24.280 19.550 24.450 19.720 ;
        RECT 25.460 19.550 25.630 19.720 ;
        RECT 25.820 19.550 25.990 19.720 ;
        RECT 26.180 19.550 26.350 19.720 ;
        RECT 26.540 19.550 26.710 19.720 ;
        RECT 26.900 19.550 27.070 19.720 ;
        RECT 27.260 19.550 27.430 19.720 ;
        RECT 27.620 19.550 27.790 19.720 ;
        RECT 27.980 19.550 28.150 19.720 ;
        RECT 28.340 19.550 28.510 19.720 ;
        RECT 29.025 19.550 29.195 19.720 ;
        RECT 29.385 19.550 29.555 19.720 ;
        RECT 29.745 19.550 29.915 19.720 ;
        RECT 30.105 19.550 30.275 19.720 ;
        RECT 30.465 19.550 30.635 19.720 ;
        RECT 30.825 19.550 30.995 19.720 ;
        RECT 31.185 19.550 31.355 19.720 ;
        RECT 31.545 19.550 31.715 19.720 ;
        RECT 31.905 19.550 32.075 19.720 ;
        RECT 32.710 19.550 32.880 19.720 ;
        RECT 33.070 19.550 33.240 19.720 ;
        RECT 33.430 19.550 33.600 19.720 ;
        RECT 33.790 19.550 33.960 19.720 ;
        RECT 34.150 19.550 34.320 19.720 ;
        RECT 34.510 19.550 34.680 19.720 ;
        RECT 34.870 19.550 35.040 19.720 ;
        RECT 35.230 19.550 35.400 19.720 ;
        RECT 35.590 19.550 35.760 19.720 ;
        RECT 36.275 19.550 36.445 19.720 ;
        RECT 36.635 19.550 36.805 19.720 ;
        RECT 36.995 19.550 37.165 19.720 ;
        RECT 37.355 19.550 37.525 19.720 ;
        RECT 37.715 19.550 37.885 19.720 ;
        RECT 38.075 19.550 38.245 19.720 ;
        RECT 38.435 19.550 38.605 19.720 ;
        RECT 38.795 19.550 38.965 19.720 ;
        RECT 39.155 19.550 39.325 19.720 ;
        RECT 40.390 19.550 40.560 19.720 ;
        RECT 40.750 19.550 40.920 19.720 ;
        RECT 41.110 19.550 41.280 19.720 ;
        RECT 41.470 19.550 41.640 19.720 ;
        RECT 41.830 19.550 42.000 19.720 ;
        RECT 42.190 19.550 42.360 19.720 ;
        RECT 42.550 19.550 42.720 19.720 ;
        RECT 42.910 19.550 43.080 19.720 ;
        RECT 43.270 19.550 43.440 19.720 ;
        RECT 43.955 19.550 44.125 19.720 ;
        RECT 44.315 19.550 44.485 19.720 ;
        RECT 44.675 19.550 44.845 19.720 ;
        RECT 45.035 19.550 45.205 19.720 ;
        RECT 45.395 19.550 45.565 19.720 ;
        RECT 45.755 19.550 45.925 19.720 ;
        RECT 46.115 19.550 46.285 19.720 ;
        RECT 46.475 19.550 46.645 19.720 ;
        RECT 46.835 19.550 47.005 19.720 ;
        RECT 47.640 19.550 47.810 19.720 ;
        RECT 48.000 19.550 48.170 19.720 ;
        RECT 48.360 19.550 48.530 19.720 ;
        RECT 48.720 19.550 48.890 19.720 ;
        RECT 49.080 19.550 49.250 19.720 ;
        RECT 49.440 19.550 49.610 19.720 ;
        RECT 49.800 19.550 49.970 19.720 ;
        RECT 50.160 19.550 50.330 19.720 ;
        RECT 50.520 19.550 50.690 19.720 ;
        RECT 51.205 19.550 51.375 19.720 ;
        RECT 51.565 19.550 51.735 19.720 ;
        RECT 51.925 19.550 52.095 19.720 ;
        RECT 52.285 19.550 52.455 19.720 ;
        RECT 52.645 19.550 52.815 19.720 ;
        RECT 53.005 19.550 53.175 19.720 ;
        RECT 53.365 19.550 53.535 19.720 ;
        RECT 53.725 19.550 53.895 19.720 ;
        RECT 54.085 19.550 54.255 19.720 ;
        RECT 55.265 19.550 55.435 19.720 ;
        RECT 55.625 19.550 55.795 19.720 ;
        RECT 55.985 19.550 56.155 19.720 ;
        RECT 56.345 19.550 56.515 19.720 ;
        RECT 56.705 19.550 56.875 19.720 ;
        RECT 57.065 19.550 57.235 19.720 ;
        RECT 57.425 19.550 57.595 19.720 ;
        RECT 57.785 19.550 57.955 19.720 ;
        RECT 58.145 19.550 58.315 19.720 ;
        RECT 58.830 19.550 59.000 19.720 ;
        RECT 59.190 19.550 59.360 19.720 ;
        RECT 59.550 19.550 59.720 19.720 ;
        RECT 59.910 19.550 60.080 19.720 ;
        RECT 60.270 19.550 60.440 19.720 ;
        RECT 60.630 19.550 60.800 19.720 ;
        RECT 60.990 19.550 61.160 19.720 ;
        RECT 61.350 19.550 61.520 19.720 ;
        RECT 61.710 19.550 61.880 19.720 ;
        RECT 62.515 19.550 62.685 19.720 ;
        RECT 62.875 19.550 63.045 19.720 ;
        RECT 63.235 19.550 63.405 19.720 ;
        RECT 63.595 19.550 63.765 19.720 ;
        RECT 63.955 19.550 64.125 19.720 ;
        RECT 64.315 19.550 64.485 19.720 ;
        RECT 64.675 19.550 64.845 19.720 ;
        RECT 65.035 19.550 65.205 19.720 ;
        RECT 65.395 19.550 65.565 19.720 ;
        RECT 66.080 19.550 66.250 19.720 ;
        RECT 66.440 19.550 66.610 19.720 ;
        RECT 66.800 19.550 66.970 19.720 ;
        RECT 67.160 19.550 67.330 19.720 ;
        RECT 67.520 19.550 67.690 19.720 ;
        RECT 67.880 19.550 68.050 19.720 ;
        RECT 68.240 19.550 68.410 19.720 ;
        RECT 68.600 19.550 68.770 19.720 ;
        RECT 68.960 19.550 69.130 19.720 ;
        RECT 70.010 19.550 70.180 19.720 ;
        RECT 70.370 19.550 70.540 19.720 ;
        RECT 70.730 19.550 70.900 19.720 ;
        RECT 71.090 19.550 71.260 19.720 ;
        RECT 71.450 19.550 71.620 19.720 ;
        RECT 71.810 19.550 71.980 19.720 ;
        RECT 72.170 19.550 72.340 19.720 ;
        RECT 72.530 19.550 72.700 19.720 ;
        RECT 72.890 19.550 73.060 19.720 ;
        RECT 73.575 19.550 73.745 19.720 ;
        RECT 73.935 19.550 74.105 19.720 ;
        RECT 74.295 19.550 74.465 19.720 ;
        RECT 74.655 19.550 74.825 19.720 ;
        RECT 75.015 19.550 75.185 19.720 ;
        RECT 75.375 19.550 75.545 19.720 ;
        RECT 75.735 19.550 75.905 19.720 ;
        RECT 76.095 19.550 76.265 19.720 ;
        RECT 76.455 19.550 76.625 19.720 ;
      LAYER met1 ;
        RECT 0.000 40.890 88.240 42.330 ;
        RECT 0.000 30.545 88.240 31.985 ;
        RECT 0.000 14.410 88.240 22.410 ;
      LAYER via ;
        RECT 75.445 41.815 75.705 42.075 ;
        RECT 75.785 41.815 76.045 42.075 ;
        RECT 76.105 41.815 76.365 42.075 ;
        RECT 76.530 41.815 76.790 42.075 ;
        RECT 76.870 41.815 77.130 42.075 ;
        RECT 75.445 41.490 75.705 41.750 ;
        RECT 75.785 41.490 76.045 41.750 ;
        RECT 76.105 41.490 76.365 41.750 ;
        RECT 76.530 41.490 76.790 41.750 ;
        RECT 76.870 41.490 77.130 41.750 ;
        RECT 75.445 41.160 75.705 41.420 ;
        RECT 75.785 41.160 76.045 41.420 ;
        RECT 76.105 41.160 76.365 41.420 ;
        RECT 76.530 41.160 76.790 41.420 ;
        RECT 76.870 41.160 77.130 41.420 ;
        RECT 75.445 31.410 75.705 31.670 ;
        RECT 75.785 31.410 76.045 31.670 ;
        RECT 76.105 31.410 76.365 31.670 ;
        RECT 76.530 31.410 76.790 31.670 ;
        RECT 76.870 31.410 77.130 31.670 ;
        RECT 75.445 31.085 75.705 31.345 ;
        RECT 75.785 31.085 76.045 31.345 ;
        RECT 76.105 31.085 76.365 31.345 ;
        RECT 76.530 31.085 76.790 31.345 ;
        RECT 76.870 31.085 77.130 31.345 ;
        RECT 75.445 30.755 75.705 31.015 ;
        RECT 75.785 30.755 76.045 31.015 ;
        RECT 76.105 30.755 76.365 31.015 ;
        RECT 76.530 30.755 76.790 31.015 ;
        RECT 76.870 30.755 77.130 31.015 ;
        RECT 75.495 21.745 75.755 22.005 ;
        RECT 75.835 21.745 76.095 22.005 ;
        RECT 76.155 21.745 76.415 22.005 ;
        RECT 76.580 21.745 76.840 22.005 ;
        RECT 76.920 21.745 77.180 22.005 ;
        RECT 75.495 21.420 75.755 21.680 ;
        RECT 75.835 21.420 76.095 21.680 ;
        RECT 76.155 21.420 76.415 21.680 ;
        RECT 76.580 21.420 76.840 21.680 ;
        RECT 76.920 21.420 77.180 21.680 ;
        RECT 75.495 21.090 75.755 21.350 ;
        RECT 75.835 21.090 76.095 21.350 ;
        RECT 76.155 21.090 76.415 21.350 ;
        RECT 76.580 21.090 76.840 21.350 ;
        RECT 76.920 21.090 77.180 21.350 ;
        RECT 75.495 20.590 75.755 20.850 ;
        RECT 75.835 20.590 76.095 20.850 ;
        RECT 76.155 20.590 76.415 20.850 ;
        RECT 76.580 20.590 76.840 20.850 ;
        RECT 76.920 20.590 77.180 20.850 ;
        RECT 75.495 20.265 75.755 20.525 ;
        RECT 75.835 20.265 76.095 20.525 ;
        RECT 76.155 20.265 76.415 20.525 ;
        RECT 76.580 20.265 76.840 20.525 ;
        RECT 76.920 20.265 77.180 20.525 ;
        RECT 75.495 19.935 75.755 20.195 ;
        RECT 75.835 19.935 76.095 20.195 ;
        RECT 76.155 19.935 76.415 20.195 ;
        RECT 76.580 19.935 76.840 20.195 ;
        RECT 76.920 19.935 77.180 20.195 ;
        RECT 75.495 19.320 75.755 19.580 ;
        RECT 75.835 19.320 76.095 19.580 ;
        RECT 76.155 19.320 76.415 19.580 ;
        RECT 76.580 19.320 76.840 19.580 ;
        RECT 76.920 19.320 77.180 19.580 ;
        RECT 75.495 18.995 75.755 19.255 ;
        RECT 75.835 18.995 76.095 19.255 ;
        RECT 76.155 18.995 76.415 19.255 ;
        RECT 76.580 18.995 76.840 19.255 ;
        RECT 76.920 18.995 77.180 19.255 ;
        RECT 75.495 18.665 75.755 18.925 ;
        RECT 75.835 18.665 76.095 18.925 ;
        RECT 76.155 18.665 76.415 18.925 ;
        RECT 76.580 18.665 76.840 18.925 ;
        RECT 76.920 18.665 77.180 18.925 ;
        RECT 75.495 18.165 75.755 18.425 ;
        RECT 75.835 18.165 76.095 18.425 ;
        RECT 76.155 18.165 76.415 18.425 ;
        RECT 76.580 18.165 76.840 18.425 ;
        RECT 76.920 18.165 77.180 18.425 ;
        RECT 75.495 17.840 75.755 18.100 ;
        RECT 75.835 17.840 76.095 18.100 ;
        RECT 76.155 17.840 76.415 18.100 ;
        RECT 76.580 17.840 76.840 18.100 ;
        RECT 76.920 17.840 77.180 18.100 ;
        RECT 75.495 17.510 75.755 17.770 ;
        RECT 75.835 17.510 76.095 17.770 ;
        RECT 76.155 17.510 76.415 17.770 ;
        RECT 76.580 17.510 76.840 17.770 ;
        RECT 76.920 17.510 77.180 17.770 ;
        RECT 75.495 16.990 75.755 17.250 ;
        RECT 75.835 16.990 76.095 17.250 ;
        RECT 76.155 16.990 76.415 17.250 ;
        RECT 76.580 16.990 76.840 17.250 ;
        RECT 76.920 16.990 77.180 17.250 ;
        RECT 75.495 16.665 75.755 16.925 ;
        RECT 75.835 16.665 76.095 16.925 ;
        RECT 76.155 16.665 76.415 16.925 ;
        RECT 76.580 16.665 76.840 16.925 ;
        RECT 76.920 16.665 77.180 16.925 ;
        RECT 75.495 16.335 75.755 16.595 ;
        RECT 75.835 16.335 76.095 16.595 ;
        RECT 76.155 16.335 76.415 16.595 ;
        RECT 76.580 16.335 76.840 16.595 ;
        RECT 76.920 16.335 77.180 16.595 ;
        RECT 75.495 15.835 75.755 16.095 ;
        RECT 75.835 15.835 76.095 16.095 ;
        RECT 76.155 15.835 76.415 16.095 ;
        RECT 76.580 15.835 76.840 16.095 ;
        RECT 76.920 15.835 77.180 16.095 ;
        RECT 75.495 15.510 75.755 15.770 ;
        RECT 75.835 15.510 76.095 15.770 ;
        RECT 76.155 15.510 76.415 15.770 ;
        RECT 76.580 15.510 76.840 15.770 ;
        RECT 76.920 15.510 77.180 15.770 ;
        RECT 75.495 15.180 75.755 15.440 ;
        RECT 75.835 15.180 76.095 15.440 ;
        RECT 76.155 15.180 76.415 15.440 ;
        RECT 76.580 15.180 76.840 15.440 ;
        RECT 76.920 15.180 77.180 15.440 ;
      LAYER met2 ;
        RECT 75.300 14.920 77.300 42.560 ;
    END
  END vdd
  PIN pad
    DIRECTION INOUT ;
    ANTENNADIFFAREA 129.675003 ;
    PORT
      LAYER li1 ;
        RECT 19.080 158.915 20.070 163.505 ;
        RECT 23.090 158.915 24.080 163.505 ;
        RECT 27.075 158.915 28.065 163.505 ;
        RECT 35.085 158.915 36.075 163.505 ;
        RECT 39.070 158.915 40.060 163.505 ;
        RECT 43.080 158.915 44.070 163.505 ;
        RECT 16.855 108.895 17.025 118.935 ;
        RECT 18.435 108.895 18.605 118.935 ;
        RECT 20.015 108.895 20.185 118.935 ;
        RECT 23.885 108.895 24.055 118.935 ;
        RECT 25.465 108.895 25.635 118.935 ;
        RECT 27.045 108.895 27.215 118.935 ;
        RECT 28.625 108.895 28.795 118.935 ;
        RECT 30.205 108.895 30.375 118.935 ;
        RECT 33.700 108.895 33.870 118.935 ;
        RECT 35.280 108.895 35.450 118.935 ;
        RECT 36.860 108.895 37.030 118.935 ;
        RECT 38.440 108.895 38.610 118.935 ;
        RECT 40.020 108.895 40.190 118.935 ;
        RECT 41.600 108.895 41.770 118.935 ;
        RECT 43.180 108.895 43.350 118.935 ;
        RECT 44.760 108.895 44.930 118.935 ;
        RECT 46.340 108.895 46.510 118.935 ;
        RECT 47.920 108.895 48.090 118.935 ;
        RECT 49.500 108.895 49.670 118.935 ;
        RECT 55.440 112.455 55.610 116.995 ;
        RECT 57.020 112.455 57.190 116.995 ;
        RECT 58.600 112.455 58.770 116.995 ;
        RECT 63.370 112.455 63.540 116.995 ;
        RECT 64.950 112.455 65.120 116.995 ;
        RECT 66.530 112.455 66.700 116.995 ;
        RECT 68.110 112.455 68.280 116.995 ;
        RECT 69.690 112.455 69.860 116.995 ;
        RECT 53.365 88.350 53.535 92.890 ;
        RECT 54.945 88.350 55.115 92.890 ;
        RECT 56.525 88.350 56.695 92.890 ;
        RECT 58.105 88.350 58.275 92.890 ;
        RECT 59.685 88.350 59.855 92.890 ;
        RECT 61.265 88.350 61.435 92.890 ;
        RECT 62.845 88.350 63.015 92.890 ;
        RECT 64.425 88.350 64.595 92.890 ;
        RECT 66.005 88.350 66.175 92.890 ;
        RECT 67.585 88.350 67.755 92.890 ;
        RECT 69.165 88.350 69.335 92.890 ;
        RECT 62.525 32.585 63.525 33.585 ;
      LAYER mcon ;
        RECT 19.280 162.930 19.450 163.100 ;
        RECT 19.705 162.930 19.875 163.100 ;
        RECT 19.280 162.570 19.450 162.740 ;
        RECT 19.705 162.570 19.875 162.740 ;
        RECT 19.280 162.210 19.450 162.380 ;
        RECT 19.705 162.210 19.875 162.380 ;
        RECT 19.280 161.850 19.450 162.020 ;
        RECT 19.705 161.850 19.875 162.020 ;
        RECT 19.280 161.490 19.450 161.660 ;
        RECT 19.705 161.490 19.875 161.660 ;
        RECT 19.280 161.130 19.450 161.300 ;
        RECT 19.705 161.130 19.875 161.300 ;
        RECT 19.280 160.770 19.450 160.940 ;
        RECT 19.705 160.770 19.875 160.940 ;
        RECT 19.280 160.410 19.450 160.580 ;
        RECT 19.705 160.410 19.875 160.580 ;
        RECT 19.280 160.050 19.450 160.220 ;
        RECT 19.705 160.050 19.875 160.220 ;
        RECT 19.280 159.690 19.450 159.860 ;
        RECT 19.705 159.690 19.875 159.860 ;
        RECT 19.280 159.330 19.450 159.500 ;
        RECT 19.705 159.330 19.875 159.500 ;
        RECT 23.310 162.930 23.480 163.100 ;
        RECT 23.735 162.930 23.905 163.100 ;
        RECT 23.310 162.570 23.480 162.740 ;
        RECT 23.735 162.570 23.905 162.740 ;
        RECT 23.310 162.210 23.480 162.380 ;
        RECT 23.735 162.210 23.905 162.380 ;
        RECT 23.310 161.850 23.480 162.020 ;
        RECT 23.735 161.850 23.905 162.020 ;
        RECT 23.310 161.490 23.480 161.660 ;
        RECT 23.735 161.490 23.905 161.660 ;
        RECT 23.310 161.130 23.480 161.300 ;
        RECT 23.735 161.130 23.905 161.300 ;
        RECT 23.310 160.770 23.480 160.940 ;
        RECT 23.735 160.770 23.905 160.940 ;
        RECT 23.310 160.410 23.480 160.580 ;
        RECT 23.735 160.410 23.905 160.580 ;
        RECT 23.310 160.050 23.480 160.220 ;
        RECT 23.735 160.050 23.905 160.220 ;
        RECT 23.310 159.690 23.480 159.860 ;
        RECT 23.735 159.690 23.905 159.860 ;
        RECT 23.310 159.330 23.480 159.500 ;
        RECT 23.735 159.330 23.905 159.500 ;
        RECT 27.275 162.930 27.445 163.100 ;
        RECT 27.700 162.930 27.870 163.100 ;
        RECT 27.275 162.570 27.445 162.740 ;
        RECT 27.700 162.570 27.870 162.740 ;
        RECT 27.275 162.210 27.445 162.380 ;
        RECT 27.700 162.210 27.870 162.380 ;
        RECT 27.275 161.850 27.445 162.020 ;
        RECT 27.700 161.850 27.870 162.020 ;
        RECT 27.275 161.490 27.445 161.660 ;
        RECT 27.700 161.490 27.870 161.660 ;
        RECT 27.275 161.130 27.445 161.300 ;
        RECT 27.700 161.130 27.870 161.300 ;
        RECT 27.275 160.770 27.445 160.940 ;
        RECT 27.700 160.770 27.870 160.940 ;
        RECT 27.275 160.410 27.445 160.580 ;
        RECT 27.700 160.410 27.870 160.580 ;
        RECT 27.275 160.050 27.445 160.220 ;
        RECT 27.700 160.050 27.870 160.220 ;
        RECT 27.275 159.690 27.445 159.860 ;
        RECT 27.700 159.690 27.870 159.860 ;
        RECT 27.275 159.330 27.445 159.500 ;
        RECT 27.700 159.330 27.870 159.500 ;
        RECT 35.280 162.930 35.450 163.100 ;
        RECT 35.705 162.930 35.875 163.100 ;
        RECT 35.280 162.570 35.450 162.740 ;
        RECT 35.705 162.570 35.875 162.740 ;
        RECT 35.280 162.210 35.450 162.380 ;
        RECT 35.705 162.210 35.875 162.380 ;
        RECT 35.280 161.850 35.450 162.020 ;
        RECT 35.705 161.850 35.875 162.020 ;
        RECT 35.280 161.490 35.450 161.660 ;
        RECT 35.705 161.490 35.875 161.660 ;
        RECT 35.280 161.130 35.450 161.300 ;
        RECT 35.705 161.130 35.875 161.300 ;
        RECT 35.280 160.770 35.450 160.940 ;
        RECT 35.705 160.770 35.875 160.940 ;
        RECT 35.280 160.410 35.450 160.580 ;
        RECT 35.705 160.410 35.875 160.580 ;
        RECT 35.280 160.050 35.450 160.220 ;
        RECT 35.705 160.050 35.875 160.220 ;
        RECT 35.280 159.690 35.450 159.860 ;
        RECT 35.705 159.690 35.875 159.860 ;
        RECT 35.280 159.330 35.450 159.500 ;
        RECT 35.705 159.330 35.875 159.500 ;
        RECT 39.245 162.930 39.415 163.100 ;
        RECT 39.670 162.930 39.840 163.100 ;
        RECT 39.245 162.570 39.415 162.740 ;
        RECT 39.670 162.570 39.840 162.740 ;
        RECT 39.245 162.210 39.415 162.380 ;
        RECT 39.670 162.210 39.840 162.380 ;
        RECT 39.245 161.850 39.415 162.020 ;
        RECT 39.670 161.850 39.840 162.020 ;
        RECT 39.245 161.490 39.415 161.660 ;
        RECT 39.670 161.490 39.840 161.660 ;
        RECT 39.245 161.130 39.415 161.300 ;
        RECT 39.670 161.130 39.840 161.300 ;
        RECT 39.245 160.770 39.415 160.940 ;
        RECT 39.670 160.770 39.840 160.940 ;
        RECT 39.245 160.410 39.415 160.580 ;
        RECT 39.670 160.410 39.840 160.580 ;
        RECT 39.245 160.050 39.415 160.220 ;
        RECT 39.670 160.050 39.840 160.220 ;
        RECT 39.245 159.690 39.415 159.860 ;
        RECT 39.670 159.690 39.840 159.860 ;
        RECT 39.245 159.330 39.415 159.500 ;
        RECT 39.670 159.330 39.840 159.500 ;
        RECT 43.275 162.930 43.445 163.100 ;
        RECT 43.700 162.930 43.870 163.100 ;
        RECT 43.275 162.570 43.445 162.740 ;
        RECT 43.700 162.570 43.870 162.740 ;
        RECT 43.275 162.210 43.445 162.380 ;
        RECT 43.700 162.210 43.870 162.380 ;
        RECT 43.275 161.850 43.445 162.020 ;
        RECT 43.700 161.850 43.870 162.020 ;
        RECT 43.275 161.490 43.445 161.660 ;
        RECT 43.700 161.490 43.870 161.660 ;
        RECT 43.275 161.130 43.445 161.300 ;
        RECT 43.700 161.130 43.870 161.300 ;
        RECT 43.275 160.770 43.445 160.940 ;
        RECT 43.700 160.770 43.870 160.940 ;
        RECT 43.275 160.410 43.445 160.580 ;
        RECT 43.700 160.410 43.870 160.580 ;
        RECT 43.275 160.050 43.445 160.220 ;
        RECT 43.700 160.050 43.870 160.220 ;
        RECT 43.275 159.690 43.445 159.860 ;
        RECT 43.700 159.690 43.870 159.860 ;
        RECT 43.275 159.330 43.445 159.500 ;
        RECT 43.700 159.330 43.870 159.500 ;
        RECT 16.855 116.610 17.025 116.780 ;
        RECT 16.855 116.250 17.025 116.420 ;
        RECT 16.855 115.890 17.025 116.060 ;
        RECT 16.855 112.670 17.025 112.840 ;
        RECT 16.855 112.310 17.025 112.480 ;
        RECT 16.855 111.950 17.025 112.120 ;
        RECT 18.435 116.610 18.605 116.780 ;
        RECT 18.435 116.250 18.605 116.420 ;
        RECT 18.435 115.890 18.605 116.060 ;
        RECT 18.435 112.670 18.605 112.840 ;
        RECT 18.435 112.310 18.605 112.480 ;
        RECT 18.435 111.950 18.605 112.120 ;
        RECT 20.015 116.610 20.185 116.780 ;
        RECT 20.015 116.250 20.185 116.420 ;
        RECT 20.015 115.890 20.185 116.060 ;
        RECT 20.015 112.670 20.185 112.840 ;
        RECT 20.015 112.310 20.185 112.480 ;
        RECT 20.015 111.950 20.185 112.120 ;
        RECT 23.885 116.610 24.055 116.780 ;
        RECT 23.885 116.250 24.055 116.420 ;
        RECT 23.885 115.890 24.055 116.060 ;
        RECT 23.885 112.670 24.055 112.840 ;
        RECT 23.885 112.310 24.055 112.480 ;
        RECT 23.885 111.950 24.055 112.120 ;
        RECT 25.465 116.610 25.635 116.780 ;
        RECT 25.465 116.250 25.635 116.420 ;
        RECT 25.465 115.890 25.635 116.060 ;
        RECT 25.465 112.670 25.635 112.840 ;
        RECT 25.465 112.310 25.635 112.480 ;
        RECT 25.465 111.950 25.635 112.120 ;
        RECT 27.045 116.610 27.215 116.780 ;
        RECT 27.045 116.250 27.215 116.420 ;
        RECT 27.045 115.890 27.215 116.060 ;
        RECT 27.045 112.670 27.215 112.840 ;
        RECT 27.045 112.310 27.215 112.480 ;
        RECT 27.045 111.950 27.215 112.120 ;
        RECT 28.625 116.610 28.795 116.780 ;
        RECT 28.625 116.250 28.795 116.420 ;
        RECT 28.625 115.890 28.795 116.060 ;
        RECT 28.625 112.670 28.795 112.840 ;
        RECT 28.625 112.310 28.795 112.480 ;
        RECT 28.625 111.950 28.795 112.120 ;
        RECT 30.205 116.610 30.375 116.780 ;
        RECT 30.205 116.250 30.375 116.420 ;
        RECT 30.205 115.890 30.375 116.060 ;
        RECT 30.205 112.670 30.375 112.840 ;
        RECT 30.205 112.310 30.375 112.480 ;
        RECT 30.205 111.950 30.375 112.120 ;
        RECT 33.700 116.610 33.870 116.780 ;
        RECT 33.700 116.250 33.870 116.420 ;
        RECT 33.700 115.890 33.870 116.060 ;
        RECT 33.700 112.670 33.870 112.840 ;
        RECT 33.700 112.310 33.870 112.480 ;
        RECT 33.700 111.950 33.870 112.120 ;
        RECT 35.280 116.610 35.450 116.780 ;
        RECT 35.280 116.250 35.450 116.420 ;
        RECT 35.280 115.890 35.450 116.060 ;
        RECT 35.280 112.670 35.450 112.840 ;
        RECT 35.280 112.310 35.450 112.480 ;
        RECT 35.280 111.950 35.450 112.120 ;
        RECT 36.860 116.610 37.030 116.780 ;
        RECT 36.860 116.250 37.030 116.420 ;
        RECT 36.860 115.890 37.030 116.060 ;
        RECT 36.860 112.670 37.030 112.840 ;
        RECT 36.860 112.310 37.030 112.480 ;
        RECT 36.860 111.950 37.030 112.120 ;
        RECT 38.440 116.610 38.610 116.780 ;
        RECT 38.440 116.250 38.610 116.420 ;
        RECT 38.440 115.890 38.610 116.060 ;
        RECT 38.440 112.670 38.610 112.840 ;
        RECT 38.440 112.310 38.610 112.480 ;
        RECT 38.440 111.950 38.610 112.120 ;
        RECT 40.020 116.610 40.190 116.780 ;
        RECT 40.020 116.250 40.190 116.420 ;
        RECT 40.020 115.890 40.190 116.060 ;
        RECT 40.020 112.670 40.190 112.840 ;
        RECT 40.020 112.310 40.190 112.480 ;
        RECT 40.020 111.950 40.190 112.120 ;
        RECT 41.600 116.610 41.770 116.780 ;
        RECT 41.600 116.250 41.770 116.420 ;
        RECT 41.600 115.890 41.770 116.060 ;
        RECT 41.600 112.670 41.770 112.840 ;
        RECT 41.600 112.310 41.770 112.480 ;
        RECT 41.600 111.950 41.770 112.120 ;
        RECT 43.180 116.610 43.350 116.780 ;
        RECT 43.180 116.250 43.350 116.420 ;
        RECT 43.180 115.890 43.350 116.060 ;
        RECT 43.180 112.670 43.350 112.840 ;
        RECT 43.180 112.310 43.350 112.480 ;
        RECT 43.180 111.950 43.350 112.120 ;
        RECT 44.760 116.610 44.930 116.780 ;
        RECT 44.760 116.250 44.930 116.420 ;
        RECT 44.760 115.890 44.930 116.060 ;
        RECT 44.760 112.670 44.930 112.840 ;
        RECT 44.760 112.310 44.930 112.480 ;
        RECT 44.760 111.950 44.930 112.120 ;
        RECT 46.340 116.610 46.510 116.780 ;
        RECT 46.340 116.250 46.510 116.420 ;
        RECT 46.340 115.890 46.510 116.060 ;
        RECT 46.340 112.670 46.510 112.840 ;
        RECT 46.340 112.310 46.510 112.480 ;
        RECT 46.340 111.950 46.510 112.120 ;
        RECT 47.920 116.610 48.090 116.780 ;
        RECT 47.920 116.250 48.090 116.420 ;
        RECT 47.920 115.890 48.090 116.060 ;
        RECT 47.920 112.670 48.090 112.840 ;
        RECT 47.920 112.310 48.090 112.480 ;
        RECT 47.920 111.950 48.090 112.120 ;
        RECT 49.500 116.610 49.670 116.780 ;
        RECT 49.500 116.250 49.670 116.420 ;
        RECT 49.500 115.890 49.670 116.060 ;
        RECT 49.500 112.670 49.670 112.840 ;
        RECT 49.500 112.310 49.670 112.480 ;
        RECT 55.440 116.620 55.610 116.790 ;
        RECT 55.440 116.260 55.610 116.430 ;
        RECT 55.440 115.900 55.610 116.070 ;
        RECT 55.440 115.540 55.610 115.710 ;
        RECT 57.020 116.620 57.190 116.790 ;
        RECT 57.020 116.260 57.190 116.430 ;
        RECT 57.020 115.900 57.190 116.070 ;
        RECT 57.020 115.540 57.190 115.710 ;
        RECT 58.600 116.620 58.770 116.790 ;
        RECT 58.600 116.260 58.770 116.430 ;
        RECT 58.600 115.900 58.770 116.070 ;
        RECT 58.600 115.540 58.770 115.710 ;
        RECT 63.370 116.620 63.540 116.790 ;
        RECT 63.370 116.260 63.540 116.430 ;
        RECT 63.370 115.900 63.540 116.070 ;
        RECT 63.370 115.540 63.540 115.710 ;
        RECT 64.950 116.620 65.120 116.790 ;
        RECT 64.950 116.260 65.120 116.430 ;
        RECT 64.950 115.900 65.120 116.070 ;
        RECT 64.950 115.540 65.120 115.710 ;
        RECT 66.530 116.620 66.700 116.790 ;
        RECT 66.530 116.260 66.700 116.430 ;
        RECT 66.530 115.900 66.700 116.070 ;
        RECT 66.530 115.540 66.700 115.710 ;
        RECT 68.110 116.620 68.280 116.790 ;
        RECT 68.110 116.260 68.280 116.430 ;
        RECT 68.110 115.900 68.280 116.070 ;
        RECT 68.110 115.540 68.280 115.710 ;
        RECT 69.690 116.620 69.860 116.790 ;
        RECT 69.690 116.260 69.860 116.430 ;
        RECT 69.690 115.900 69.860 116.070 ;
        RECT 69.690 115.540 69.860 115.710 ;
        RECT 49.500 111.950 49.670 112.120 ;
        RECT 53.365 89.635 53.535 89.805 ;
        RECT 53.365 89.275 53.535 89.445 ;
        RECT 53.365 88.915 53.535 89.085 ;
        RECT 53.365 88.555 53.535 88.725 ;
        RECT 54.945 89.635 55.115 89.805 ;
        RECT 54.945 89.275 55.115 89.445 ;
        RECT 54.945 88.915 55.115 89.085 ;
        RECT 54.945 88.555 55.115 88.725 ;
        RECT 56.525 89.635 56.695 89.805 ;
        RECT 56.525 89.275 56.695 89.445 ;
        RECT 56.525 88.915 56.695 89.085 ;
        RECT 56.525 88.555 56.695 88.725 ;
        RECT 58.105 89.635 58.275 89.805 ;
        RECT 58.105 89.275 58.275 89.445 ;
        RECT 58.105 88.915 58.275 89.085 ;
        RECT 58.105 88.555 58.275 88.725 ;
        RECT 59.685 89.635 59.855 89.805 ;
        RECT 59.685 89.275 59.855 89.445 ;
        RECT 59.685 88.915 59.855 89.085 ;
        RECT 59.685 88.555 59.855 88.725 ;
        RECT 61.265 89.635 61.435 89.805 ;
        RECT 61.265 89.275 61.435 89.445 ;
        RECT 61.265 88.915 61.435 89.085 ;
        RECT 61.265 88.555 61.435 88.725 ;
        RECT 62.845 89.635 63.015 89.805 ;
        RECT 62.845 89.275 63.015 89.445 ;
        RECT 62.845 88.915 63.015 89.085 ;
        RECT 62.845 88.555 63.015 88.725 ;
        RECT 64.425 89.635 64.595 89.805 ;
        RECT 64.425 89.275 64.595 89.445 ;
        RECT 64.425 88.915 64.595 89.085 ;
        RECT 64.425 88.555 64.595 88.725 ;
        RECT 66.005 89.635 66.175 89.805 ;
        RECT 66.005 89.275 66.175 89.445 ;
        RECT 66.005 88.915 66.175 89.085 ;
        RECT 66.005 88.555 66.175 88.725 ;
        RECT 67.585 89.635 67.755 89.805 ;
        RECT 67.585 89.275 67.755 89.445 ;
        RECT 67.585 88.915 67.755 89.085 ;
        RECT 67.585 88.555 67.755 88.725 ;
        RECT 69.165 89.635 69.335 89.805 ;
        RECT 69.165 89.275 69.335 89.445 ;
        RECT 69.165 88.915 69.335 89.085 ;
        RECT 69.165 88.555 69.335 88.725 ;
        RECT 62.740 33.160 62.910 33.330 ;
        RECT 63.210 33.160 63.380 33.330 ;
        RECT 62.740 32.800 62.910 32.970 ;
        RECT 63.210 32.800 63.380 32.970 ;
      LAYER met1 ;
        RECT 19.020 159.115 20.145 163.255 ;
        RECT 23.055 159.155 24.180 163.305 ;
        RECT 26.995 159.125 28.050 163.255 ;
        RECT 35.100 159.125 36.155 163.255 ;
        RECT 38.970 159.155 40.095 163.305 ;
        RECT 43.005 159.115 44.130 163.255 ;
        RECT 11.175 115.665 71.120 116.975 ;
        RECT 55.165 115.230 59.015 115.665 ;
        RECT 63.265 115.230 69.990 115.665 ;
        RECT 11.175 111.725 49.890 113.035 ;
        RECT 53.335 88.370 69.430 90.115 ;
        RECT 62.515 32.465 63.590 33.595 ;
      LAYER via ;
        RECT 19.295 162.470 19.555 162.730 ;
        RECT 19.635 162.470 19.895 162.730 ;
        RECT 19.295 162.145 19.555 162.405 ;
        RECT 19.635 162.145 19.895 162.405 ;
        RECT 19.295 161.815 19.555 162.075 ;
        RECT 19.635 161.815 19.895 162.075 ;
        RECT 19.295 161.325 19.555 161.585 ;
        RECT 19.635 161.325 19.895 161.585 ;
        RECT 19.295 161.000 19.555 161.260 ;
        RECT 19.635 161.000 19.895 161.260 ;
        RECT 19.295 160.670 19.555 160.930 ;
        RECT 19.635 160.670 19.895 160.930 ;
        RECT 19.295 160.165 19.555 160.425 ;
        RECT 19.635 160.165 19.895 160.425 ;
        RECT 19.295 159.840 19.555 160.100 ;
        RECT 19.635 159.840 19.895 160.100 ;
        RECT 19.295 159.510 19.555 159.770 ;
        RECT 19.635 159.510 19.895 159.770 ;
        RECT 23.355 162.470 23.615 162.730 ;
        RECT 23.695 162.470 23.955 162.730 ;
        RECT 23.355 162.145 23.615 162.405 ;
        RECT 23.695 162.145 23.955 162.405 ;
        RECT 23.355 161.815 23.615 162.075 ;
        RECT 23.695 161.815 23.955 162.075 ;
        RECT 23.355 161.325 23.615 161.585 ;
        RECT 23.695 161.325 23.955 161.585 ;
        RECT 23.355 161.000 23.615 161.260 ;
        RECT 23.695 161.000 23.955 161.260 ;
        RECT 23.355 160.670 23.615 160.930 ;
        RECT 23.695 160.670 23.955 160.930 ;
        RECT 23.355 160.165 23.615 160.425 ;
        RECT 23.695 160.165 23.955 160.425 ;
        RECT 23.355 159.840 23.615 160.100 ;
        RECT 23.695 159.840 23.955 160.100 ;
        RECT 23.355 159.510 23.615 159.770 ;
        RECT 23.695 159.510 23.955 159.770 ;
        RECT 27.230 162.470 27.490 162.730 ;
        RECT 27.570 162.470 27.830 162.730 ;
        RECT 27.230 162.145 27.490 162.405 ;
        RECT 27.570 162.145 27.830 162.405 ;
        RECT 27.230 161.815 27.490 162.075 ;
        RECT 27.570 161.815 27.830 162.075 ;
        RECT 27.230 161.325 27.490 161.585 ;
        RECT 27.570 161.325 27.830 161.585 ;
        RECT 27.230 161.000 27.490 161.260 ;
        RECT 27.570 161.000 27.830 161.260 ;
        RECT 27.230 160.670 27.490 160.930 ;
        RECT 27.570 160.670 27.830 160.930 ;
        RECT 27.230 160.165 27.490 160.425 ;
        RECT 27.570 160.165 27.830 160.425 ;
        RECT 27.230 159.840 27.490 160.100 ;
        RECT 27.570 159.840 27.830 160.100 ;
        RECT 27.230 159.510 27.490 159.770 ;
        RECT 27.570 159.510 27.830 159.770 ;
        RECT 35.315 162.470 35.575 162.730 ;
        RECT 35.655 162.470 35.915 162.730 ;
        RECT 35.315 162.145 35.575 162.405 ;
        RECT 35.655 162.145 35.915 162.405 ;
        RECT 35.315 161.815 35.575 162.075 ;
        RECT 35.655 161.815 35.915 162.075 ;
        RECT 35.315 161.325 35.575 161.585 ;
        RECT 35.655 161.325 35.915 161.585 ;
        RECT 35.315 161.000 35.575 161.260 ;
        RECT 35.655 161.000 35.915 161.260 ;
        RECT 35.315 160.670 35.575 160.930 ;
        RECT 35.655 160.670 35.915 160.930 ;
        RECT 35.315 160.165 35.575 160.425 ;
        RECT 35.655 160.165 35.915 160.425 ;
        RECT 35.315 159.840 35.575 160.100 ;
        RECT 35.655 159.840 35.915 160.100 ;
        RECT 35.315 159.510 35.575 159.770 ;
        RECT 35.655 159.510 35.915 159.770 ;
        RECT 39.375 162.470 39.635 162.730 ;
        RECT 39.715 162.470 39.975 162.730 ;
        RECT 39.375 162.145 39.635 162.405 ;
        RECT 39.715 162.145 39.975 162.405 ;
        RECT 39.375 161.815 39.635 162.075 ;
        RECT 39.715 161.815 39.975 162.075 ;
        RECT 39.375 161.325 39.635 161.585 ;
        RECT 39.715 161.325 39.975 161.585 ;
        RECT 39.375 161.000 39.635 161.260 ;
        RECT 39.715 161.000 39.975 161.260 ;
        RECT 39.375 160.670 39.635 160.930 ;
        RECT 39.715 160.670 39.975 160.930 ;
        RECT 39.375 160.165 39.635 160.425 ;
        RECT 39.715 160.165 39.975 160.425 ;
        RECT 39.375 159.840 39.635 160.100 ;
        RECT 39.715 159.840 39.975 160.100 ;
        RECT 39.375 159.510 39.635 159.770 ;
        RECT 39.715 159.510 39.975 159.770 ;
        RECT 43.250 162.470 43.510 162.730 ;
        RECT 43.590 162.470 43.850 162.730 ;
        RECT 43.250 162.145 43.510 162.405 ;
        RECT 43.590 162.145 43.850 162.405 ;
        RECT 43.250 161.815 43.510 162.075 ;
        RECT 43.590 161.815 43.850 162.075 ;
        RECT 43.250 161.325 43.510 161.585 ;
        RECT 43.590 161.325 43.850 161.585 ;
        RECT 43.250 161.000 43.510 161.260 ;
        RECT 43.590 161.000 43.850 161.260 ;
        RECT 43.250 160.670 43.510 160.930 ;
        RECT 43.590 160.670 43.850 160.930 ;
        RECT 43.250 160.165 43.510 160.425 ;
        RECT 43.590 160.165 43.850 160.425 ;
        RECT 43.250 159.840 43.510 160.100 ;
        RECT 43.590 159.840 43.850 160.100 ;
        RECT 43.250 159.510 43.510 159.770 ;
        RECT 43.590 159.510 43.850 159.770 ;
        RECT 17.995 116.140 18.255 116.400 ;
        RECT 18.335 116.140 18.595 116.400 ;
        RECT 18.655 116.140 18.915 116.400 ;
        RECT 19.060 116.140 19.320 116.400 ;
        RECT 19.400 116.140 19.660 116.400 ;
        RECT 19.720 116.140 19.980 116.400 ;
        RECT 26.240 116.180 26.500 116.440 ;
        RECT 26.580 116.180 26.840 116.440 ;
        RECT 26.900 116.180 27.160 116.440 ;
        RECT 27.305 116.180 27.565 116.440 ;
        RECT 27.645 116.180 27.905 116.440 ;
        RECT 27.965 116.180 28.225 116.440 ;
        RECT 28.450 116.180 28.710 116.440 ;
        RECT 28.790 116.180 29.050 116.440 ;
        RECT 36.360 116.305 36.620 116.565 ;
        RECT 36.700 116.305 36.960 116.565 ;
        RECT 37.020 116.305 37.280 116.565 ;
        RECT 37.425 116.305 37.685 116.565 ;
        RECT 37.765 116.305 38.025 116.565 ;
        RECT 38.085 116.305 38.345 116.565 ;
        RECT 38.570 116.305 38.830 116.565 ;
        RECT 38.910 116.305 39.170 116.565 ;
        RECT 41.715 116.545 41.975 116.805 ;
        RECT 42.055 116.545 42.315 116.805 ;
        RECT 42.375 116.545 42.635 116.805 ;
        RECT 42.780 116.545 43.040 116.805 ;
        RECT 43.120 116.545 43.380 116.805 ;
        RECT 43.440 116.545 43.700 116.805 ;
        RECT 43.925 116.545 44.185 116.805 ;
        RECT 44.265 116.545 44.525 116.805 ;
        RECT 44.585 116.545 44.845 116.805 ;
        RECT 44.990 116.545 45.250 116.805 ;
        RECT 45.330 116.545 45.590 116.805 ;
        RECT 46.020 116.545 46.280 116.805 ;
        RECT 46.360 116.545 46.620 116.805 ;
        RECT 46.680 116.545 46.940 116.805 ;
        RECT 47.085 116.545 47.345 116.805 ;
        RECT 47.425 116.545 47.685 116.805 ;
        RECT 47.745 116.545 48.005 116.805 ;
        RECT 48.230 116.545 48.490 116.805 ;
        RECT 48.570 116.545 48.830 116.805 ;
        RECT 48.890 116.545 49.150 116.805 ;
        RECT 49.295 116.545 49.555 116.805 ;
        RECT 49.635 116.545 49.895 116.805 ;
        RECT 41.715 116.220 41.975 116.480 ;
        RECT 42.055 116.220 42.315 116.480 ;
        RECT 42.375 116.220 42.635 116.480 ;
        RECT 42.780 116.220 43.040 116.480 ;
        RECT 43.120 116.220 43.380 116.480 ;
        RECT 43.440 116.220 43.700 116.480 ;
        RECT 43.925 116.220 44.185 116.480 ;
        RECT 44.265 116.220 44.525 116.480 ;
        RECT 44.585 116.220 44.845 116.480 ;
        RECT 44.990 116.220 45.250 116.480 ;
        RECT 45.330 116.220 45.590 116.480 ;
        RECT 46.020 116.220 46.280 116.480 ;
        RECT 46.360 116.220 46.620 116.480 ;
        RECT 46.680 116.220 46.940 116.480 ;
        RECT 47.085 116.220 47.345 116.480 ;
        RECT 47.425 116.220 47.685 116.480 ;
        RECT 47.745 116.220 48.005 116.480 ;
        RECT 48.230 116.220 48.490 116.480 ;
        RECT 48.570 116.220 48.830 116.480 ;
        RECT 48.890 116.220 49.150 116.480 ;
        RECT 49.295 116.220 49.555 116.480 ;
        RECT 49.635 116.220 49.895 116.480 ;
        RECT 41.715 115.890 41.975 116.150 ;
        RECT 42.055 115.890 42.315 116.150 ;
        RECT 42.375 115.890 42.635 116.150 ;
        RECT 42.780 115.890 43.040 116.150 ;
        RECT 43.120 115.890 43.380 116.150 ;
        RECT 43.440 115.890 43.700 116.150 ;
        RECT 43.925 115.890 44.185 116.150 ;
        RECT 44.265 115.890 44.525 116.150 ;
        RECT 44.585 115.890 44.845 116.150 ;
        RECT 44.990 115.890 45.250 116.150 ;
        RECT 45.330 115.890 45.590 116.150 ;
        RECT 46.020 115.890 46.280 116.150 ;
        RECT 46.360 115.890 46.620 116.150 ;
        RECT 46.680 115.890 46.940 116.150 ;
        RECT 47.085 115.890 47.345 116.150 ;
        RECT 47.425 115.890 47.685 116.150 ;
        RECT 47.745 115.890 48.005 116.150 ;
        RECT 48.230 115.890 48.490 116.150 ;
        RECT 48.570 115.890 48.830 116.150 ;
        RECT 48.890 115.890 49.150 116.150 ;
        RECT 49.295 115.890 49.555 116.150 ;
        RECT 49.635 115.890 49.895 116.150 ;
        RECT 17.995 112.240 18.255 112.500 ;
        RECT 18.335 112.240 18.595 112.500 ;
        RECT 18.655 112.240 18.915 112.500 ;
        RECT 19.060 112.240 19.320 112.500 ;
        RECT 19.400 112.240 19.660 112.500 ;
        RECT 19.720 112.240 19.980 112.500 ;
        RECT 26.240 112.235 26.500 112.495 ;
        RECT 26.580 112.235 26.840 112.495 ;
        RECT 26.900 112.235 27.160 112.495 ;
        RECT 27.305 112.235 27.565 112.495 ;
        RECT 27.645 112.235 27.905 112.495 ;
        RECT 27.965 112.235 28.225 112.495 ;
        RECT 28.450 112.235 28.710 112.495 ;
        RECT 28.790 112.235 29.050 112.495 ;
        RECT 36.360 112.180 36.620 112.440 ;
        RECT 36.700 112.180 36.960 112.440 ;
        RECT 37.020 112.180 37.280 112.440 ;
        RECT 37.425 112.180 37.685 112.440 ;
        RECT 37.765 112.180 38.025 112.440 ;
        RECT 38.085 112.180 38.345 112.440 ;
        RECT 38.570 112.180 38.830 112.440 ;
        RECT 38.910 112.180 39.170 112.440 ;
        RECT 55.335 89.640 55.595 89.900 ;
        RECT 55.675 89.640 55.935 89.900 ;
        RECT 56.240 89.640 56.500 89.900 ;
        RECT 56.580 89.640 56.840 89.900 ;
        RECT 56.900 89.640 57.160 89.900 ;
        RECT 57.305 89.640 57.565 89.900 ;
        RECT 57.645 89.640 57.905 89.900 ;
        RECT 57.965 89.640 58.225 89.900 ;
        RECT 58.450 89.640 58.710 89.900 ;
        RECT 55.335 89.315 55.595 89.575 ;
        RECT 55.675 89.315 55.935 89.575 ;
        RECT 56.240 89.315 56.500 89.575 ;
        RECT 56.580 89.315 56.840 89.575 ;
        RECT 56.900 89.315 57.160 89.575 ;
        RECT 57.305 89.315 57.565 89.575 ;
        RECT 57.645 89.315 57.905 89.575 ;
        RECT 57.965 89.315 58.225 89.575 ;
        RECT 58.450 89.315 58.710 89.575 ;
        RECT 55.335 88.890 55.595 89.150 ;
        RECT 55.675 88.890 55.935 89.150 ;
        RECT 56.240 88.890 56.500 89.150 ;
        RECT 56.580 88.890 56.840 89.150 ;
        RECT 56.900 88.890 57.160 89.150 ;
        RECT 57.305 88.890 57.565 89.150 ;
        RECT 57.645 88.890 57.905 89.150 ;
        RECT 57.965 88.890 58.225 89.150 ;
        RECT 58.450 88.890 58.710 89.150 ;
        RECT 55.335 88.565 55.595 88.825 ;
        RECT 55.675 88.565 55.935 88.825 ;
        RECT 56.240 88.565 56.500 88.825 ;
        RECT 56.580 88.565 56.840 88.825 ;
        RECT 56.900 88.565 57.160 88.825 ;
        RECT 57.305 88.565 57.565 88.825 ;
        RECT 57.645 88.565 57.905 88.825 ;
        RECT 57.965 88.565 58.225 88.825 ;
        RECT 58.450 88.565 58.710 88.825 ;
        RECT 62.740 33.285 63.000 33.545 ;
        RECT 63.070 33.285 63.330 33.545 ;
        RECT 62.740 32.945 63.000 33.205 ;
        RECT 63.070 32.945 63.330 33.205 ;
        RECT 62.740 32.625 63.000 32.885 ;
        RECT 63.070 32.625 63.330 32.885 ;
      LAYER met2 ;
        RECT 28.375 162.970 34.375 182.520 ;
        RECT 19.130 159.330 44.295 162.970 ;
        RECT 29.000 152.885 33.000 159.330 ;
        RECT 29.000 148.885 45.265 152.885 ;
        RECT 41.265 122.800 45.265 148.885 ;
        RECT 41.265 120.800 60.500 122.800 ;
        RECT 41.265 118.405 45.265 120.800 ;
        RECT 17.775 116.005 20.960 116.505 ;
        RECT 25.830 116.050 29.380 116.550 ;
        RECT 36.150 116.175 39.250 116.675 ;
        RECT 17.775 112.645 18.275 116.005 ;
        RECT 17.775 112.145 20.195 112.645 ;
        RECT 25.830 112.640 26.330 116.050 ;
        RECT 25.830 112.140 29.205 112.640 ;
        RECT 36.150 112.565 36.650 116.175 ;
        RECT 41.265 114.405 50.595 118.405 ;
        RECT 36.150 112.065 40.510 112.565 ;
        RECT 58.500 90.230 60.500 120.800 ;
        RECT 54.710 88.230 60.500 90.230 ;
        RECT 56.480 52.590 56.820 88.230 ;
        RECT 56.480 52.250 64.750 52.590 ;
        RECT 62.195 33.240 63.670 33.845 ;
        RECT 64.410 33.240 64.750 52.250 ;
        RECT 62.195 32.900 64.750 33.240 ;
        RECT 62.195 32.235 63.670 32.900 ;
    END
  END pad
  PIN in
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.040000 ;
    PORT
      LAYER li1 ;
        RECT 56.180 28.275 56.590 31.240 ;
        RECT 57.820 28.275 58.150 31.240 ;
        RECT 59.380 28.275 59.710 31.240 ;
        RECT 60.940 28.275 61.270 31.240 ;
        RECT 62.500 28.275 62.830 31.240 ;
        RECT 64.060 28.275 64.390 31.240 ;
        RECT 65.620 28.275 65.950 31.240 ;
        RECT 67.180 28.275 67.510 31.240 ;
      LAYER mcon ;
        RECT 56.340 29.805 56.510 29.975 ;
        RECT 57.900 29.805 58.070 29.975 ;
        RECT 59.460 29.805 59.630 29.975 ;
        RECT 61.020 29.805 61.190 29.975 ;
        RECT 62.580 29.805 62.750 29.975 ;
        RECT 64.140 29.805 64.310 29.975 ;
        RECT 65.700 29.805 65.870 29.975 ;
        RECT 67.260 29.805 67.430 29.975 ;
      LAYER met1 ;
        RECT 56.280 29.975 56.570 30.005 ;
        RECT 57.840 29.975 58.130 30.005 ;
        RECT 59.400 29.975 59.690 30.005 ;
        RECT 60.960 29.975 61.250 30.005 ;
        RECT 62.520 29.975 62.810 30.005 ;
        RECT 63.335 29.975 67.505 30.075 ;
        RECT 56.280 29.805 67.505 29.975 ;
        RECT 56.280 29.775 56.570 29.805 ;
        RECT 57.840 29.775 58.130 29.805 ;
        RECT 59.400 29.775 59.690 29.805 ;
        RECT 60.960 29.775 61.250 29.805 ;
        RECT 62.520 29.775 62.810 29.805 ;
        RECT 63.335 29.720 67.505 29.805 ;
      LAYER via ;
        RECT 63.810 29.755 64.070 30.015 ;
        RECT 64.150 29.755 64.410 30.015 ;
        RECT 64.470 29.755 64.730 30.015 ;
        RECT 64.980 29.755 65.240 30.015 ;
        RECT 65.320 29.755 65.580 30.015 ;
        RECT 65.640 29.755 65.900 30.015 ;
      LAYER met2 ;
        RECT 63.275 29.730 67.455 30.070 ;
        RECT 67.115 0.000 67.455 29.730 ;
    END
  END in
  PIN oe_l
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.960000 ;
    PORT
      LAYER li1 ;
        RECT 15.410 39.485 16.850 39.735 ;
        RECT 40.250 39.485 41.690 39.735 ;
        RECT 61.640 39.485 63.080 39.735 ;
        RECT 25.775 29.140 29.080 29.390 ;
      LAYER mcon ;
        RECT 15.650 39.500 15.820 39.670 ;
        RECT 16.010 39.500 16.180 39.670 ;
        RECT 16.370 39.500 16.540 39.670 ;
        RECT 40.335 39.530 40.505 39.700 ;
        RECT 40.705 39.530 40.875 39.700 ;
        RECT 41.065 39.530 41.235 39.700 ;
        RECT 41.425 39.530 41.595 39.700 ;
        RECT 61.735 39.530 61.905 39.700 ;
        RECT 62.105 39.530 62.275 39.700 ;
        RECT 62.465 39.530 62.635 39.700 ;
        RECT 62.825 39.530 62.995 39.700 ;
        RECT 27.830 29.175 28.000 29.345 ;
        RECT 28.190 29.175 28.360 29.345 ;
      LAYER met1 ;
        RECT 15.375 39.055 16.940 39.755 ;
        RECT 40.230 39.055 41.795 39.755 ;
        RECT 61.630 39.055 63.195 39.755 ;
        RECT 8.730 35.155 74.215 35.655 ;
        RECT 27.600 29.120 29.165 29.410 ;
        RECT 8.730 24.860 74.215 25.360 ;
      LAYER via ;
        RECT 15.535 39.135 15.795 39.395 ;
        RECT 15.875 39.135 16.135 39.395 ;
        RECT 16.195 39.135 16.455 39.395 ;
        RECT 16.535 39.135 16.795 39.395 ;
        RECT 41.050 39.135 41.310 39.395 ;
        RECT 41.390 39.135 41.650 39.395 ;
        RECT 61.790 39.135 62.050 39.395 ;
        RECT 62.130 39.135 62.390 39.395 ;
        RECT 9.060 35.290 9.320 35.550 ;
        RECT 9.400 35.290 9.660 35.550 ;
        RECT 9.720 35.290 9.980 35.550 ;
        RECT 15.565 35.290 15.825 35.550 ;
        RECT 15.905 35.290 16.165 35.550 ;
        RECT 16.225 35.290 16.485 35.550 ;
        RECT 16.565 35.290 16.825 35.550 ;
        RECT 41.080 35.290 41.340 35.550 ;
        RECT 41.420 35.290 41.680 35.550 ;
        RECT 61.820 35.290 62.080 35.550 ;
        RECT 62.160 35.290 62.420 35.550 ;
        RECT 27.825 29.130 28.085 29.390 ;
        RECT 28.165 29.130 28.425 29.390 ;
        RECT 9.060 24.985 9.320 25.245 ;
        RECT 9.400 24.985 9.660 25.245 ;
        RECT 9.720 24.985 9.980 25.245 ;
        RECT 27.855 24.945 28.115 25.205 ;
        RECT 28.195 24.945 28.455 25.205 ;
      LAYER met2 ;
        RECT 9.010 0.000 10.010 35.910 ;
        RECT 15.395 35.110 16.875 39.510 ;
        RECT 40.920 35.110 41.730 39.510 ;
        RECT 61.650 35.110 62.575 39.510 ;
        RECT 27.700 24.765 28.615 29.585 ;
    END
  END oe_l
  PIN out_l
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.940000 ;
    PORT
      LAYER li1 ;
        RECT 17.735 39.485 19.355 39.735 ;
        RECT 31.995 39.485 33.615 39.735 ;
        RECT 50.855 39.485 52.475 39.735 ;
        RECT 21.570 29.140 23.230 29.340 ;
        RECT 38.130 29.140 39.790 29.340 ;
        RECT 52.390 29.140 54.050 29.340 ;
      LAYER mcon ;
        RECT 17.980 39.500 18.150 39.670 ;
        RECT 18.340 39.500 18.510 39.670 ;
        RECT 18.700 39.500 18.870 39.670 ;
        RECT 19.070 39.500 19.240 39.670 ;
        RECT 32.180 39.530 32.350 39.700 ;
        RECT 32.550 39.530 32.720 39.700 ;
        RECT 32.910 39.530 33.080 39.700 ;
        RECT 33.270 39.530 33.440 39.700 ;
        RECT 51.040 39.525 51.210 39.695 ;
        RECT 51.410 39.525 51.580 39.695 ;
        RECT 51.770 39.525 51.940 39.695 ;
        RECT 52.130 39.525 52.300 39.695 ;
        RECT 22.390 29.155 22.560 29.325 ;
        RECT 22.750 29.155 22.920 29.325 ;
        RECT 38.670 29.160 38.840 29.330 ;
        RECT 39.030 29.160 39.200 29.330 ;
        RECT 39.390 29.160 39.560 29.330 ;
        RECT 52.580 29.155 52.750 29.325 ;
        RECT 52.940 29.155 53.110 29.325 ;
        RECT 53.310 29.155 53.480 29.325 ;
      LAYER met1 ;
        RECT 17.825 39.055 19.390 39.755 ;
        RECT 31.960 39.055 33.625 39.755 ;
        RECT 50.820 39.055 52.485 39.755 ;
        RECT 8.730 34.155 74.215 34.655 ;
        RECT 21.665 29.095 23.145 29.385 ;
        RECT 38.385 28.710 39.855 29.410 ;
        RECT 52.365 28.710 54.030 29.410 ;
        RECT 8.730 23.860 74.215 24.360 ;
      LAYER via ;
        RECT 17.985 39.135 18.245 39.395 ;
        RECT 18.325 39.135 18.585 39.395 ;
        RECT 18.645 39.135 18.905 39.395 ;
        RECT 18.985 39.135 19.245 39.395 ;
        RECT 32.220 39.135 32.480 39.395 ;
        RECT 32.560 39.135 32.820 39.395 ;
        RECT 32.880 39.135 33.140 39.395 ;
        RECT 33.220 39.135 33.480 39.395 ;
        RECT 51.080 39.135 51.340 39.395 ;
        RECT 51.420 39.135 51.680 39.395 ;
        RECT 51.740 39.135 52.000 39.395 ;
        RECT 52.080 39.135 52.340 39.395 ;
        RECT 10.820 34.290 11.080 34.550 ;
        RECT 11.160 34.290 11.420 34.550 ;
        RECT 11.480 34.290 11.740 34.550 ;
        RECT 18.015 34.265 18.275 34.525 ;
        RECT 18.355 34.265 18.615 34.525 ;
        RECT 18.675 34.265 18.935 34.525 ;
        RECT 19.015 34.265 19.275 34.525 ;
        RECT 32.250 34.285 32.510 34.545 ;
        RECT 32.590 34.285 32.850 34.545 ;
        RECT 32.910 34.285 33.170 34.545 ;
        RECT 33.250 34.285 33.510 34.545 ;
        RECT 51.110 34.285 51.370 34.545 ;
        RECT 51.450 34.285 51.710 34.545 ;
        RECT 51.770 34.285 52.030 34.545 ;
        RECT 52.110 34.285 52.370 34.545 ;
        RECT 22.350 29.105 22.610 29.365 ;
        RECT 22.690 29.105 22.950 29.365 ;
        RECT 38.435 28.790 38.695 29.050 ;
        RECT 38.775 28.790 39.035 29.050 ;
        RECT 39.095 28.790 39.355 29.050 ;
        RECT 39.435 28.790 39.695 29.050 ;
        RECT 52.510 28.790 52.770 29.050 ;
        RECT 52.850 28.790 53.110 29.050 ;
        RECT 53.170 28.790 53.430 29.050 ;
        RECT 53.510 28.790 53.770 29.050 ;
        RECT 10.820 23.985 11.080 24.245 ;
        RECT 11.160 23.985 11.420 24.245 ;
        RECT 11.480 23.985 11.740 24.245 ;
        RECT 22.350 23.930 22.610 24.190 ;
        RECT 22.690 23.930 22.950 24.190 ;
        RECT 38.405 23.940 38.665 24.200 ;
        RECT 38.745 23.940 39.005 24.200 ;
        RECT 39.065 23.940 39.325 24.200 ;
        RECT 39.405 23.940 39.665 24.200 ;
        RECT 52.480 23.940 52.740 24.200 ;
        RECT 52.820 23.940 53.080 24.200 ;
        RECT 53.140 23.940 53.400 24.200 ;
        RECT 53.480 23.940 53.740 24.200 ;
      LAYER met2 ;
        RECT 10.770 0.000 11.770 34.905 ;
        RECT 17.845 34.085 19.325 39.510 ;
        RECT 32.080 34.105 33.560 39.510 ;
        RECT 50.940 34.105 52.420 39.510 ;
        RECT 22.155 23.680 23.025 29.585 ;
        RECT 38.355 23.760 39.835 29.165 ;
        RECT 52.430 23.760 53.910 29.165 ;
    END
  END out_l
  PIN strong_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 59.135 39.485 60.755 39.735 ;
      LAYER mcon ;
        RECT 59.285 39.530 59.455 39.700 ;
        RECT 59.655 39.530 59.825 39.700 ;
        RECT 60.015 39.530 60.185 39.700 ;
        RECT 60.375 39.530 60.545 39.700 ;
      LAYER met1 ;
        RECT 59.220 39.055 60.785 39.755 ;
      LAYER via ;
        RECT 59.380 39.135 59.640 39.395 ;
        RECT 59.720 39.135 59.980 39.395 ;
        RECT 60.040 39.135 60.300 39.395 ;
        RECT 60.380 39.135 60.640 39.395 ;
      LAYER met2 ;
        RECT 59.240 0.000 60.720 39.510 ;
    END
  END strong_enable
  PIN med_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 42.575 39.485 44.195 39.735 ;
      LAYER mcon ;
        RECT 42.735 39.530 42.905 39.700 ;
        RECT 43.105 39.530 43.275 39.700 ;
        RECT 43.465 39.530 43.635 39.700 ;
        RECT 43.825 39.530 43.995 39.700 ;
      LAYER met1 ;
        RECT 42.670 39.055 44.235 39.755 ;
      LAYER via ;
        RECT 42.830 39.135 43.090 39.395 ;
        RECT 43.170 39.135 43.430 39.395 ;
        RECT 43.490 39.135 43.750 39.395 ;
        RECT 43.830 39.135 44.090 39.395 ;
      LAYER met2 ;
        RECT 42.690 0.000 44.170 39.510 ;
    END
  END med_enable
  OBS
      LAYER pwell ;
        RECT 15.590 38.515 19.460 39.425 ;
        RECT 21.360 38.515 23.550 39.425 ;
        RECT 27.800 38.515 29.990 39.425 ;
        RECT 31.890 38.515 35.760 39.425 ;
        RECT 36.080 38.515 38.270 39.425 ;
        RECT 40.430 38.515 44.300 39.425 ;
        RECT 46.660 38.515 48.850 39.425 ;
        RECT 50.750 38.515 54.620 39.425 ;
        RECT 54.940 38.515 57.130 39.425 ;
        RECT 59.030 38.515 62.900 39.425 ;
        RECT 19.145 38.325 19.315 38.515 ;
        RECT 21.020 38.350 21.130 38.470 ;
        RECT 21.450 38.325 21.620 38.515 ;
        RECT 25.160 38.350 25.270 38.470 ;
        RECT 27.460 38.350 27.570 38.470 ;
        RECT 29.730 38.325 29.900 38.515 ;
        RECT 31.600 38.350 31.710 38.470 ;
        RECT 32.035 38.325 32.205 38.515 ;
        RECT 38.010 38.325 38.180 38.515 ;
        RECT 39.880 38.350 39.990 38.470 ;
        RECT 43.985 38.325 44.155 38.515 ;
        RECT 46.320 38.350 46.430 38.470 ;
        RECT 48.590 38.325 48.760 38.515 ;
        RECT 50.460 38.350 50.570 38.470 ;
        RECT 50.895 38.325 51.065 38.515 ;
        RECT 56.870 38.325 57.040 38.515 ;
        RECT 58.740 38.350 58.850 38.470 ;
        RECT 59.175 38.325 59.345 38.515 ;
        RECT 15.145 28.170 17.335 29.080 ;
        RECT 19.475 28.170 23.365 29.080 ;
        RECT 25.265 28.170 27.455 29.080 ;
        RECT 31.705 28.170 33.895 29.080 ;
        RECT 36.035 28.170 39.925 29.080 ;
        RECT 45.965 28.170 48.155 29.080 ;
        RECT 50.295 28.170 54.185 29.080 ;
        RECT 14.805 28.005 14.915 28.125 ;
        RECT 17.075 27.980 17.245 28.170 ;
        RECT 18.945 28.005 19.055 28.125 ;
        RECT 23.050 27.980 23.220 28.170 ;
        RECT 24.925 28.005 25.035 28.125 ;
        RECT 27.195 27.980 27.365 28.170 ;
        RECT 29.065 28.005 29.175 28.125 ;
        RECT 29.985 28.005 30.095 28.125 ;
        RECT 33.635 27.980 33.805 28.170 ;
        RECT 34.125 28.005 34.235 28.125 ;
        RECT 39.610 27.980 39.780 28.170 ;
        RECT 40.565 28.005 40.675 28.125 ;
        RECT 42.405 28.005 42.515 28.125 ;
        RECT 44.245 28.005 44.355 28.125 ;
        RECT 47.895 27.980 48.065 28.170 ;
        RECT 48.385 28.005 48.495 28.125 ;
        RECT 53.870 27.980 54.040 28.170 ;
      LAYER li1 ;
        RECT 16.295 119.150 16.795 120.605 ;
        RECT 17.085 119.150 17.585 120.605 ;
        RECT 17.875 119.150 18.375 120.605 ;
        RECT 18.665 119.150 19.165 120.605 ;
        RECT 19.455 119.150 19.955 120.605 ;
        RECT 20.245 119.150 20.745 120.605 ;
        RECT 23.325 119.150 23.825 120.605 ;
        RECT 24.115 119.150 24.615 120.605 ;
        RECT 24.905 119.150 25.405 120.605 ;
        RECT 25.695 119.150 26.195 120.605 ;
        RECT 26.485 119.150 26.985 120.605 ;
        RECT 27.275 119.150 27.775 120.605 ;
        RECT 28.065 119.150 28.565 120.605 ;
        RECT 28.855 119.150 29.355 120.605 ;
        RECT 29.645 119.150 30.145 120.605 ;
        RECT 33.140 119.150 33.640 120.605 ;
        RECT 33.930 119.150 34.430 120.605 ;
        RECT 34.720 119.150 35.220 120.605 ;
        RECT 35.510 119.150 36.010 120.605 ;
        RECT 36.300 119.150 36.800 120.605 ;
        RECT 37.090 119.150 37.590 120.605 ;
        RECT 37.880 119.150 38.380 120.605 ;
        RECT 38.670 119.150 39.170 120.605 ;
        RECT 39.460 119.150 39.960 120.605 ;
        RECT 40.250 119.150 40.750 120.605 ;
        RECT 41.040 119.150 41.540 120.605 ;
        RECT 41.830 119.150 42.330 120.605 ;
        RECT 42.620 119.150 43.120 120.605 ;
        RECT 43.410 119.150 43.910 120.605 ;
        RECT 44.200 119.150 44.700 120.605 ;
        RECT 44.990 119.150 45.490 120.605 ;
        RECT 45.780 119.150 46.280 120.605 ;
        RECT 46.570 119.150 47.070 120.605 ;
        RECT 47.360 119.150 47.860 120.605 ;
        RECT 48.150 119.150 48.650 120.605 ;
        RECT 48.940 119.150 49.440 120.605 ;
        RECT 49.730 119.150 50.230 120.605 ;
        RECT 54.880 117.165 59.330 118.700 ;
        RECT 62.810 117.165 69.630 118.700 ;
        RECT 54.880 110.735 59.330 112.285 ;
        RECT 62.810 110.735 69.630 112.285 ;
        RECT 16.295 107.560 16.795 108.680 ;
        RECT 17.085 107.560 17.585 108.680 ;
        RECT 17.875 107.560 18.375 108.680 ;
        RECT 18.665 107.560 19.165 108.680 ;
        RECT 19.455 107.560 19.955 108.680 ;
        RECT 20.245 107.560 20.745 108.680 ;
        RECT 23.325 107.560 23.825 108.680 ;
        RECT 24.115 107.560 24.615 108.680 ;
        RECT 24.905 107.560 25.405 108.680 ;
        RECT 25.695 107.560 26.195 108.680 ;
        RECT 26.485 107.560 26.985 108.680 ;
        RECT 27.275 107.560 27.775 108.680 ;
        RECT 28.065 107.560 28.565 108.680 ;
        RECT 28.855 107.560 29.355 108.680 ;
        RECT 29.645 107.560 30.145 108.680 ;
        RECT 33.140 107.560 33.640 108.680 ;
        RECT 33.930 107.560 34.430 108.680 ;
        RECT 34.720 107.560 35.220 108.680 ;
        RECT 35.510 107.560 36.010 108.680 ;
        RECT 36.300 107.560 36.800 108.680 ;
        RECT 37.090 107.560 37.590 108.680 ;
        RECT 37.880 107.560 38.380 108.680 ;
        RECT 38.670 107.560 39.170 108.680 ;
        RECT 39.460 107.560 39.960 108.680 ;
        RECT 40.250 107.560 40.750 108.680 ;
        RECT 41.040 107.560 41.540 108.680 ;
        RECT 41.830 107.560 42.330 108.680 ;
        RECT 42.620 107.560 43.120 108.680 ;
        RECT 43.410 107.560 43.910 108.680 ;
        RECT 44.200 107.560 44.700 108.680 ;
        RECT 44.990 107.560 45.490 108.680 ;
        RECT 45.780 107.560 46.280 108.680 ;
        RECT 46.570 107.560 47.070 108.680 ;
        RECT 47.360 107.560 47.860 108.680 ;
        RECT 48.150 107.560 48.650 108.680 ;
        RECT 48.940 107.560 49.440 108.680 ;
        RECT 49.730 107.560 50.230 108.680 ;
        RECT 16.375 104.095 16.705 105.750 ;
        RECT 18.015 104.095 18.265 105.750 ;
        RECT 16.375 103.925 19.050 104.095 ;
        RECT 15.460 103.575 18.170 103.745 ;
        RECT 18.350 103.545 19.050 103.925 ;
        RECT 18.350 103.395 18.520 103.545 ;
        RECT 16.375 103.225 18.520 103.395 ;
        RECT 16.375 102.490 16.625 103.225 ;
        RECT 17.935 102.490 18.520 103.225 ;
        RECT 20.075 102.790 20.405 105.750 ;
        RECT 20.575 103.560 21.465 103.890 ;
        RECT 21.635 102.790 21.965 105.750 ;
        RECT 22.135 103.560 23.025 103.890 ;
        RECT 23.195 102.790 23.525 105.750 ;
        RECT 23.695 103.560 24.585 103.890 ;
        RECT 24.755 102.790 25.085 105.750 ;
        RECT 25.255 103.560 26.145 103.890 ;
        RECT 26.315 102.790 26.645 105.750 ;
        RECT 26.815 103.560 27.705 103.890 ;
        RECT 27.875 102.790 28.205 105.750 ;
        RECT 28.375 103.560 29.265 103.890 ;
        RECT 29.435 102.790 29.765 105.750 ;
        RECT 29.935 103.560 30.825 103.890 ;
        RECT 30.995 102.790 31.325 105.750 ;
        RECT 33.655 104.095 33.985 105.750 ;
        RECT 35.295 104.095 35.545 105.750 ;
        RECT 33.655 103.925 36.330 104.095 ;
        RECT 32.740 103.575 35.450 103.745 ;
        RECT 35.630 103.545 36.330 103.925 ;
        RECT 35.630 103.395 35.800 103.545 ;
        RECT 33.655 103.225 35.800 103.395 ;
        RECT 33.655 102.490 33.905 103.225 ;
        RECT 35.215 102.490 35.800 103.225 ;
        RECT 37.355 102.790 37.685 105.750 ;
        RECT 37.855 103.560 38.745 103.890 ;
        RECT 38.915 102.790 39.245 105.750 ;
        RECT 39.415 103.560 40.305 103.890 ;
        RECT 40.475 102.790 40.805 105.750 ;
        RECT 40.975 103.560 41.865 103.890 ;
        RECT 42.035 102.790 42.365 105.750 ;
        RECT 42.535 103.560 43.425 103.890 ;
        RECT 43.595 102.790 43.925 105.750 ;
        RECT 44.095 103.560 44.985 103.890 ;
        RECT 45.155 102.790 45.485 105.750 ;
        RECT 45.655 103.560 46.545 103.890 ;
        RECT 46.715 102.790 47.045 105.750 ;
        RECT 47.215 103.560 48.105 103.890 ;
        RECT 48.275 102.790 48.605 105.750 ;
        RECT 50.935 104.095 51.265 105.750 ;
        RECT 52.575 104.095 52.825 105.750 ;
        RECT 50.935 103.925 53.610 104.095 ;
        RECT 50.020 103.575 52.730 103.745 ;
        RECT 52.910 103.545 53.610 103.925 ;
        RECT 52.910 103.395 53.080 103.545 ;
        RECT 50.935 103.225 53.080 103.395 ;
        RECT 50.935 102.490 51.185 103.225 ;
        RECT 52.495 102.490 53.080 103.225 ;
        RECT 54.635 102.790 54.965 105.750 ;
        RECT 55.135 103.560 56.025 103.890 ;
        RECT 56.195 102.790 56.525 105.750 ;
        RECT 56.695 103.560 57.585 103.890 ;
        RECT 57.755 102.790 58.085 105.750 ;
        RECT 58.255 103.560 59.145 103.890 ;
        RECT 59.315 102.790 59.645 105.750 ;
        RECT 59.815 103.560 60.705 103.890 ;
        RECT 60.875 102.790 61.205 105.750 ;
        RECT 61.375 103.560 62.265 103.890 ;
        RECT 62.435 102.790 62.765 105.750 ;
        RECT 62.935 103.560 63.825 103.890 ;
        RECT 63.995 102.790 64.325 105.750 ;
        RECT 64.495 103.560 65.385 103.890 ;
        RECT 65.555 102.790 65.885 105.750 ;
        RECT 16.375 100.765 16.625 101.500 ;
        RECT 17.935 100.765 18.520 101.500 ;
        RECT 16.375 100.595 18.520 100.765 ;
        RECT 18.350 100.445 18.520 100.595 ;
        RECT 15.460 100.245 18.170 100.415 ;
        RECT 18.350 100.065 19.050 100.445 ;
        RECT 16.375 99.895 19.050 100.065 ;
        RECT 16.375 98.240 16.705 99.895 ;
        RECT 18.015 98.240 18.265 99.895 ;
        RECT 20.075 98.240 20.405 101.200 ;
        RECT 20.575 100.100 21.465 100.430 ;
        RECT 21.635 98.240 21.965 101.200 ;
        RECT 22.135 100.100 23.025 100.430 ;
        RECT 23.195 98.240 23.525 101.200 ;
        RECT 23.695 100.100 24.585 100.430 ;
        RECT 24.755 98.240 25.085 101.200 ;
        RECT 25.255 100.100 26.145 100.430 ;
        RECT 26.315 98.240 26.645 101.200 ;
        RECT 26.815 100.100 27.705 100.430 ;
        RECT 27.875 98.240 28.205 101.200 ;
        RECT 28.375 100.100 29.265 100.430 ;
        RECT 29.435 98.240 29.765 101.200 ;
        RECT 29.935 100.100 30.825 100.430 ;
        RECT 30.995 98.240 31.325 101.200 ;
        RECT 33.655 100.765 33.905 101.500 ;
        RECT 35.215 100.765 35.800 101.500 ;
        RECT 33.655 100.595 35.800 100.765 ;
        RECT 35.630 100.445 35.800 100.595 ;
        RECT 32.740 100.245 35.450 100.415 ;
        RECT 35.630 100.065 36.330 100.445 ;
        RECT 33.655 99.895 36.330 100.065 ;
        RECT 33.655 98.240 33.985 99.895 ;
        RECT 35.295 98.240 35.545 99.895 ;
        RECT 37.355 98.240 37.685 101.200 ;
        RECT 37.855 100.100 38.745 100.430 ;
        RECT 38.915 98.240 39.245 101.200 ;
        RECT 39.415 100.100 40.305 100.430 ;
        RECT 40.475 98.240 40.805 101.200 ;
        RECT 40.975 100.100 41.865 100.430 ;
        RECT 42.035 98.240 42.365 101.200 ;
        RECT 42.535 100.100 43.425 100.430 ;
        RECT 43.595 98.240 43.925 101.200 ;
        RECT 44.095 100.100 44.985 100.430 ;
        RECT 45.155 98.240 45.485 101.200 ;
        RECT 45.655 100.100 46.545 100.430 ;
        RECT 46.715 98.240 47.045 101.200 ;
        RECT 47.215 100.100 48.105 100.430 ;
        RECT 48.275 98.240 48.605 101.200 ;
        RECT 50.935 100.765 51.185 101.500 ;
        RECT 52.495 100.765 53.080 101.500 ;
        RECT 50.935 100.595 53.080 100.765 ;
        RECT 52.910 100.445 53.080 100.595 ;
        RECT 50.020 100.245 52.730 100.415 ;
        RECT 52.910 100.065 53.610 100.445 ;
        RECT 50.935 99.895 53.610 100.065 ;
        RECT 50.935 98.240 51.265 99.895 ;
        RECT 52.575 98.240 52.825 99.895 ;
        RECT 54.635 98.240 54.965 101.200 ;
        RECT 55.135 100.100 56.025 100.430 ;
        RECT 56.195 98.240 56.525 101.200 ;
        RECT 56.695 100.100 57.585 100.430 ;
        RECT 57.755 98.240 58.085 101.200 ;
        RECT 58.255 100.100 59.145 100.430 ;
        RECT 59.315 98.240 59.645 101.200 ;
        RECT 59.815 100.100 60.705 100.430 ;
        RECT 60.875 98.240 61.205 101.200 ;
        RECT 61.375 100.100 62.265 100.430 ;
        RECT 62.435 98.240 62.765 101.200 ;
        RECT 62.935 100.100 63.825 100.430 ;
        RECT 63.995 98.240 64.325 101.200 ;
        RECT 64.495 100.100 65.385 100.430 ;
        RECT 65.555 98.240 65.885 101.200 ;
        RECT 16.755 95.720 17.735 96.220 ;
        RECT 19.210 95.720 20.220 96.220 ;
        RECT 22.515 95.720 23.495 96.220 ;
        RECT 24.970 95.720 25.980 96.220 ;
        RECT 28.275 95.720 29.255 96.220 ;
        RECT 30.730 95.720 31.740 96.220 ;
        RECT 34.035 95.720 35.015 96.220 ;
        RECT 36.490 95.720 37.500 96.220 ;
        RECT 39.795 95.720 40.775 96.220 ;
        RECT 42.250 95.720 43.260 96.220 ;
        RECT 45.555 95.720 46.535 96.220 ;
        RECT 48.010 95.720 49.020 96.220 ;
        RECT 16.755 94.930 17.735 95.430 ;
        RECT 19.210 94.930 20.230 95.430 ;
        RECT 22.515 94.930 23.495 95.430 ;
        RECT 24.970 94.930 25.990 95.430 ;
        RECT 28.275 94.930 29.255 95.430 ;
        RECT 30.730 94.930 31.750 95.430 ;
        RECT 34.035 94.930 35.015 95.430 ;
        RECT 36.490 94.930 37.510 95.430 ;
        RECT 39.795 94.930 40.775 95.430 ;
        RECT 42.250 94.930 43.270 95.430 ;
        RECT 45.555 94.930 46.535 95.430 ;
        RECT 48.010 94.930 49.030 95.430 ;
        RECT 17.955 94.700 18.995 94.870 ;
        RECT 23.715 94.700 24.755 94.870 ;
        RECT 29.475 94.700 30.515 94.870 ;
        RECT 35.235 94.700 36.275 94.870 ;
        RECT 40.995 94.700 42.035 94.870 ;
        RECT 46.755 94.700 47.795 94.870 ;
        RECT 16.530 93.430 20.220 93.700 ;
        RECT 22.290 93.430 25.980 93.700 ;
        RECT 28.050 93.430 31.740 93.700 ;
        RECT 33.810 93.430 37.500 93.700 ;
        RECT 39.570 93.430 43.260 93.700 ;
        RECT 45.330 93.430 49.020 93.700 ;
        RECT 52.805 93.060 69.105 94.610 ;
        RECT 17.895 92.145 18.935 92.315 ;
        RECT 23.655 92.145 24.695 92.315 ;
        RECT 29.415 92.145 30.455 92.315 ;
        RECT 35.175 92.145 36.215 92.315 ;
        RECT 40.935 92.145 41.975 92.315 ;
        RECT 46.695 92.145 47.735 92.315 ;
        RECT 16.655 91.585 17.725 92.085 ;
        RECT 19.105 91.585 20.195 92.085 ;
        RECT 22.415 91.585 23.485 92.085 ;
        RECT 24.865 91.585 25.955 92.085 ;
        RECT 28.175 91.585 29.245 92.085 ;
        RECT 30.625 91.585 31.715 92.085 ;
        RECT 33.935 91.585 35.005 92.085 ;
        RECT 36.385 91.585 37.475 92.085 ;
        RECT 39.695 91.585 40.765 92.085 ;
        RECT 42.145 91.585 43.235 92.085 ;
        RECT 45.455 91.585 46.525 92.085 ;
        RECT 47.905 91.585 48.995 92.085 ;
        RECT 16.655 90.505 17.725 91.005 ;
        RECT 19.105 90.505 20.115 91.005 ;
        RECT 22.415 90.505 23.485 91.005 ;
        RECT 24.865 90.505 25.875 91.005 ;
        RECT 28.175 90.505 29.245 91.005 ;
        RECT 30.625 90.505 31.635 91.005 ;
        RECT 33.935 90.505 35.005 91.005 ;
        RECT 36.385 90.505 37.395 91.005 ;
        RECT 39.695 90.505 40.765 91.005 ;
        RECT 42.145 90.505 43.155 91.005 ;
        RECT 45.455 90.505 46.525 91.005 ;
        RECT 47.905 90.505 48.915 91.005 ;
        RECT 17.895 90.275 18.935 90.445 ;
        RECT 23.655 90.275 24.695 90.445 ;
        RECT 29.415 90.275 30.455 90.445 ;
        RECT 35.175 90.275 36.215 90.445 ;
        RECT 40.935 90.275 41.975 90.445 ;
        RECT 46.695 90.275 47.735 90.445 ;
        RECT 16.530 88.960 20.220 89.230 ;
        RECT 22.290 88.960 25.980 89.230 ;
        RECT 28.050 88.960 31.740 89.230 ;
        RECT 33.810 88.960 37.500 89.230 ;
        RECT 39.570 88.960 43.260 89.230 ;
        RECT 45.330 88.960 49.020 89.230 ;
        RECT 17.955 87.535 18.995 87.705 ;
        RECT 23.715 87.535 24.755 87.705 ;
        RECT 29.475 87.535 30.515 87.705 ;
        RECT 35.235 87.535 36.275 87.705 ;
        RECT 40.995 87.535 42.035 87.705 ;
        RECT 46.755 87.535 47.795 87.705 ;
        RECT 16.655 86.975 17.735 87.475 ;
        RECT 19.210 86.975 20.220 87.475 ;
        RECT 22.415 86.975 23.495 87.475 ;
        RECT 24.970 86.975 25.980 87.475 ;
        RECT 28.175 86.975 29.255 87.475 ;
        RECT 30.730 86.975 31.740 87.475 ;
        RECT 33.935 86.975 35.015 87.475 ;
        RECT 36.490 86.975 37.500 87.475 ;
        RECT 39.695 86.975 40.775 87.475 ;
        RECT 42.250 86.975 43.260 87.475 ;
        RECT 45.455 86.975 46.535 87.475 ;
        RECT 48.010 86.975 49.020 87.475 ;
        RECT 52.805 86.645 69.105 88.180 ;
        RECT 16.655 85.895 17.735 86.395 ;
        RECT 19.210 85.895 20.220 86.395 ;
        RECT 22.415 85.895 23.495 86.395 ;
        RECT 24.970 85.895 25.980 86.395 ;
        RECT 28.175 85.895 29.255 86.395 ;
        RECT 30.730 85.895 31.740 86.395 ;
        RECT 33.935 85.895 35.015 86.395 ;
        RECT 36.490 85.895 37.500 86.395 ;
        RECT 39.695 85.895 40.775 86.395 ;
        RECT 42.250 85.895 43.260 86.395 ;
        RECT 45.455 85.895 46.535 86.395 ;
        RECT 48.010 85.895 49.020 86.395 ;
        RECT 16.100 40.075 16.430 40.875 ;
        RECT 16.940 40.075 17.270 40.875 ;
        RECT 17.780 40.075 18.110 40.875 ;
        RECT 18.620 40.075 18.950 40.875 ;
        RECT 16.100 39.905 18.950 40.075 ;
        RECT 17.020 39.485 17.555 39.905 ;
        RECT 19.715 39.735 21.070 40.585 ;
        RECT 21.870 40.075 22.200 40.875 ;
        RECT 22.710 40.095 23.040 40.875 ;
        RECT 26.170 40.095 27.460 40.490 ;
        RECT 28.310 40.095 28.640 40.875 ;
        RECT 22.710 40.075 24.985 40.095 ;
        RECT 21.870 39.905 24.985 40.075 ;
        RECT 19.715 39.485 23.040 39.735 ;
        RECT 15.680 38.875 15.930 39.295 ;
        RECT 17.020 39.215 17.270 39.485 ;
        RECT 23.210 39.315 24.985 39.905 ;
        RECT 16.100 39.045 17.270 39.215 ;
        RECT 17.440 39.125 19.375 39.315 ;
        RECT 17.440 38.875 17.690 39.125 ;
        RECT 15.680 38.665 17.690 38.875 ;
        RECT 18.200 38.665 18.530 39.125 ;
        RECT 19.040 38.665 19.375 39.125 ;
        RECT 21.870 39.135 24.985 39.315 ;
        RECT 26.170 40.075 28.640 40.095 ;
        RECT 29.150 40.075 29.480 40.875 ;
        RECT 26.170 39.905 29.480 40.075 ;
        RECT 26.170 39.315 28.140 39.905 ;
        RECT 30.225 39.735 31.650 40.575 ;
        RECT 32.400 40.075 32.730 40.875 ;
        RECT 33.240 40.075 33.570 40.875 ;
        RECT 34.080 40.075 34.410 40.875 ;
        RECT 34.920 40.075 35.250 40.875 ;
        RECT 36.590 40.095 36.920 40.875 ;
        RECT 32.400 39.905 35.250 40.075 ;
        RECT 36.155 40.075 36.920 40.095 ;
        RECT 37.430 40.075 37.760 40.875 ;
        RECT 36.155 39.905 37.760 40.075 ;
        RECT 28.310 39.485 31.650 39.735 ;
        RECT 33.795 39.485 34.330 39.905 ;
        RECT 36.155 39.735 36.420 39.905 ;
        RECT 38.535 39.735 39.860 40.505 ;
        RECT 40.940 40.075 41.270 40.875 ;
        RECT 41.780 40.075 42.110 40.875 ;
        RECT 42.620 40.075 42.950 40.875 ;
        RECT 43.460 40.075 43.790 40.875 ;
        RECT 40.940 39.905 43.790 40.075 ;
        RECT 45.030 40.095 46.320 40.490 ;
        RECT 47.170 40.095 47.500 40.875 ;
        RECT 45.030 40.075 47.500 40.095 ;
        RECT 48.010 40.075 48.340 40.875 ;
        RECT 45.030 39.905 48.340 40.075 ;
        RECT 34.500 39.485 36.420 39.735 ;
        RECT 36.590 39.485 39.860 39.735 ;
        RECT 41.860 39.485 42.395 39.905 ;
        RECT 30.225 39.335 31.650 39.485 ;
        RECT 26.170 39.135 29.480 39.315 ;
        RECT 21.870 38.665 22.200 39.135 ;
        RECT 22.710 38.665 23.040 39.135 ;
        RECT 28.310 38.665 28.640 39.135 ;
        RECT 29.150 38.665 29.480 39.135 ;
        RECT 31.975 39.125 33.910 39.315 ;
        RECT 31.975 38.665 32.310 39.125 ;
        RECT 32.820 38.665 33.150 39.125 ;
        RECT 33.660 38.875 33.910 39.125 ;
        RECT 34.080 39.215 34.330 39.485 ;
        RECT 36.155 39.315 36.420 39.485 ;
        RECT 34.080 39.045 35.250 39.215 ;
        RECT 35.420 38.875 35.670 39.295 ;
        RECT 36.155 39.135 37.760 39.315 ;
        RECT 33.660 38.665 35.670 38.875 ;
        RECT 36.590 38.665 36.920 39.135 ;
        RECT 37.430 38.665 37.760 39.135 ;
        RECT 40.520 38.875 40.770 39.295 ;
        RECT 41.860 39.215 42.110 39.485 ;
        RECT 45.030 39.315 47.000 39.905 ;
        RECT 49.085 39.735 50.510 40.575 ;
        RECT 51.260 40.075 51.590 40.875 ;
        RECT 52.100 40.075 52.430 40.875 ;
        RECT 52.940 40.075 53.270 40.875 ;
        RECT 53.780 40.075 54.110 40.875 ;
        RECT 55.450 40.095 55.780 40.875 ;
        RECT 51.260 39.905 54.110 40.075 ;
        RECT 55.015 40.075 55.780 40.095 ;
        RECT 56.290 40.075 56.620 40.875 ;
        RECT 55.015 39.905 56.620 40.075 ;
        RECT 47.170 39.485 50.510 39.735 ;
        RECT 52.655 39.485 53.190 39.905 ;
        RECT 55.015 39.735 55.280 39.905 ;
        RECT 57.395 39.735 58.720 40.505 ;
        RECT 59.540 40.075 59.870 40.875 ;
        RECT 60.380 40.075 60.710 40.875 ;
        RECT 61.220 40.075 61.550 40.875 ;
        RECT 62.060 40.075 62.390 40.875 ;
        RECT 59.540 39.905 62.390 40.075 ;
        RECT 53.360 39.485 55.280 39.735 ;
        RECT 55.450 39.485 58.720 39.735 ;
        RECT 60.935 39.485 61.470 39.905 ;
        RECT 49.085 39.335 50.510 39.485 ;
        RECT 40.940 39.045 42.110 39.215 ;
        RECT 42.280 39.125 44.215 39.315 ;
        RECT 45.030 39.135 48.340 39.315 ;
        RECT 42.280 38.875 42.530 39.125 ;
        RECT 40.520 38.665 42.530 38.875 ;
        RECT 43.040 38.665 43.370 39.125 ;
        RECT 43.880 38.665 44.215 39.125 ;
        RECT 47.170 38.665 47.500 39.135 ;
        RECT 48.010 38.665 48.340 39.135 ;
        RECT 50.835 39.125 52.770 39.315 ;
        RECT 50.835 38.665 51.170 39.125 ;
        RECT 51.680 38.665 52.010 39.125 ;
        RECT 52.520 38.875 52.770 39.125 ;
        RECT 52.940 39.215 53.190 39.485 ;
        RECT 55.015 39.315 55.280 39.485 ;
        RECT 52.940 39.045 54.110 39.215 ;
        RECT 54.280 38.875 54.530 39.295 ;
        RECT 55.015 39.135 56.620 39.315 ;
        RECT 52.520 38.665 54.530 38.875 ;
        RECT 55.450 38.665 55.780 39.135 ;
        RECT 56.290 38.665 56.620 39.135 ;
        RECT 59.115 39.125 61.050 39.315 ;
        RECT 59.115 38.665 59.450 39.125 ;
        RECT 59.960 38.665 60.290 39.125 ;
        RECT 60.800 38.875 61.050 39.125 ;
        RECT 61.220 39.215 61.470 39.485 ;
        RECT 61.220 39.045 62.390 39.215 ;
        RECT 62.560 38.875 62.810 39.295 ;
        RECT 60.800 38.665 62.810 38.875 ;
        RECT 73.525 32.585 74.505 33.585 ;
        RECT 15.655 29.750 15.985 30.530 ;
        RECT 13.710 29.730 15.985 29.750 ;
        RECT 16.495 29.730 16.825 30.530 ;
        RECT 19.480 30.360 21.575 30.530 ;
        RECT 19.480 29.980 19.895 30.360 ;
        RECT 20.065 29.810 20.235 30.190 ;
        RECT 20.405 30.000 20.735 30.360 ;
        RECT 20.905 29.810 21.075 30.190 ;
        RECT 13.710 29.560 16.825 29.730 ;
        RECT 13.710 28.970 15.485 29.560 ;
        RECT 17.805 29.510 21.075 29.810 ;
        RECT 21.245 29.730 21.575 30.360 ;
        RECT 22.165 29.730 22.335 30.530 ;
        RECT 23.005 29.730 23.280 30.530 ;
        RECT 25.775 29.750 26.105 30.530 ;
        RECT 21.245 29.520 23.280 29.730 ;
        RECT 23.635 29.730 26.105 29.750 ;
        RECT 26.615 29.730 26.945 30.530 ;
        RECT 23.635 29.560 26.945 29.730 ;
        RECT 17.805 29.390 19.715 29.510 ;
        RECT 15.655 29.140 19.715 29.390 ;
        RECT 19.885 29.140 21.250 29.340 ;
        RECT 17.805 28.970 19.715 29.140 ;
        RECT 23.635 28.970 25.605 29.560 ;
        RECT 30.120 29.390 31.445 30.160 ;
        RECT 32.215 29.750 32.545 30.530 ;
        RECT 31.780 29.730 32.545 29.750 ;
        RECT 33.055 29.730 33.385 30.530 ;
        RECT 36.040 30.360 38.135 30.530 ;
        RECT 31.780 29.560 33.385 29.730 ;
        RECT 34.255 29.810 35.580 30.160 ;
        RECT 36.040 29.980 36.455 30.360 ;
        RECT 36.625 29.810 36.795 30.190 ;
        RECT 36.965 30.000 37.295 30.360 ;
        RECT 37.465 29.810 37.635 30.190 ;
        RECT 31.780 29.390 32.045 29.560 ;
        RECT 34.255 29.510 37.635 29.810 ;
        RECT 37.805 29.730 38.135 30.360 ;
        RECT 38.725 29.730 38.895 30.530 ;
        RECT 39.565 29.730 39.840 30.530 ;
        RECT 37.805 29.520 39.840 29.730 ;
        RECT 34.255 29.390 36.275 29.510 ;
        RECT 30.120 29.140 32.045 29.390 ;
        RECT 32.215 29.140 36.275 29.390 ;
        RECT 44.380 29.390 45.705 30.160 ;
        RECT 46.475 29.750 46.805 30.530 ;
        RECT 46.040 29.730 46.805 29.750 ;
        RECT 47.315 29.730 47.645 30.530 ;
        RECT 50.300 30.360 52.395 30.530 ;
        RECT 46.040 29.560 47.645 29.730 ;
        RECT 48.515 29.810 49.840 30.160 ;
        RECT 50.300 29.980 50.715 30.360 ;
        RECT 50.885 29.810 51.055 30.190 ;
        RECT 51.225 30.000 51.555 30.360 ;
        RECT 51.725 29.810 51.895 30.190 ;
        RECT 46.040 29.390 46.305 29.560 ;
        RECT 48.515 29.510 51.895 29.810 ;
        RECT 52.065 29.730 52.395 30.360 ;
        RECT 52.985 29.730 53.155 30.530 ;
        RECT 53.825 29.730 54.100 30.530 ;
        RECT 68.790 29.750 69.140 31.240 ;
        RECT 70.370 29.750 70.680 31.240 ;
        RECT 71.920 29.750 72.230 31.240 ;
        RECT 52.065 29.520 54.100 29.730 ;
        RECT 48.515 29.390 50.535 29.510 ;
        RECT 36.445 29.140 37.810 29.340 ;
        RECT 44.380 29.140 46.305 29.390 ;
        RECT 46.475 29.140 50.535 29.390 ;
        RECT 67.730 29.470 72.230 29.750 ;
        RECT 50.705 29.140 52.070 29.340 ;
        RECT 31.780 28.970 32.045 29.140 ;
        RECT 34.255 28.970 36.275 29.140 ;
        RECT 46.040 28.970 46.305 29.140 ;
        RECT 48.515 28.970 50.535 29.140 ;
        RECT 56.890 29.050 57.560 29.380 ;
        RECT 58.450 29.050 59.120 29.380 ;
        RECT 60.010 29.050 60.680 29.380 ;
        RECT 61.570 29.050 62.240 29.380 ;
        RECT 63.130 29.050 63.800 29.380 ;
        RECT 64.690 29.050 65.360 29.380 ;
        RECT 66.250 29.050 66.920 29.380 ;
        RECT 13.710 28.790 16.825 28.970 ;
        RECT 17.805 28.790 22.835 28.970 ;
        RECT 23.635 28.790 26.945 28.970 ;
        RECT 31.780 28.790 33.385 28.970 ;
        RECT 34.255 28.790 39.395 28.970 ;
        RECT 46.040 28.790 47.645 28.970 ;
        RECT 48.515 28.790 53.655 28.970 ;
        RECT 15.655 28.320 15.985 28.790 ;
        RECT 16.495 28.320 16.825 28.790 ;
        RECT 19.985 28.320 20.315 28.790 ;
        RECT 20.825 28.320 21.155 28.790 ;
        RECT 21.665 28.320 21.995 28.790 ;
        RECT 22.505 28.320 22.835 28.790 ;
        RECT 25.775 28.320 26.105 28.790 ;
        RECT 26.615 28.320 26.945 28.790 ;
        RECT 32.215 28.320 32.545 28.790 ;
        RECT 33.055 28.320 33.385 28.790 ;
        RECT 36.545 28.320 36.875 28.790 ;
        RECT 37.385 28.320 37.715 28.790 ;
        RECT 38.225 28.320 38.555 28.790 ;
        RECT 39.065 28.320 39.395 28.790 ;
        RECT 46.475 28.320 46.805 28.790 ;
        RECT 47.315 28.320 47.645 28.790 ;
        RECT 50.805 28.320 51.135 28.790 ;
        RECT 51.645 28.320 51.975 28.790 ;
        RECT 52.485 28.320 52.815 28.790 ;
        RECT 53.325 28.320 53.655 28.790 ;
        RECT 67.730 28.895 68.280 29.470 ;
        RECT 68.450 29.065 72.860 29.300 ;
        RECT 67.730 28.680 72.265 28.895 ;
        RECT 68.810 28.215 69.055 28.680 ;
        RECT 70.290 28.215 70.680 28.680 ;
        RECT 71.910 28.240 72.265 28.680 ;
      LAYER mcon ;
        RECT 16.460 120.315 16.630 120.485 ;
        RECT 16.460 119.950 16.630 120.120 ;
        RECT 16.460 119.540 16.630 119.710 ;
        RECT 17.250 120.315 17.420 120.485 ;
        RECT 17.250 119.950 17.420 120.120 ;
        RECT 17.250 119.540 17.420 119.710 ;
        RECT 18.040 120.315 18.210 120.485 ;
        RECT 18.040 119.950 18.210 120.120 ;
        RECT 18.040 119.540 18.210 119.710 ;
        RECT 18.830 120.315 19.000 120.485 ;
        RECT 18.830 119.950 19.000 120.120 ;
        RECT 18.830 119.540 19.000 119.710 ;
        RECT 19.620 120.315 19.790 120.485 ;
        RECT 19.620 119.950 19.790 120.120 ;
        RECT 19.620 119.540 19.790 119.710 ;
        RECT 20.410 120.315 20.580 120.485 ;
        RECT 20.410 119.950 20.580 120.120 ;
        RECT 20.410 119.540 20.580 119.710 ;
        RECT 23.490 120.315 23.660 120.485 ;
        RECT 23.490 119.950 23.660 120.120 ;
        RECT 23.490 119.540 23.660 119.710 ;
        RECT 24.280 120.315 24.450 120.485 ;
        RECT 24.280 119.950 24.450 120.120 ;
        RECT 24.280 119.540 24.450 119.710 ;
        RECT 25.070 120.315 25.240 120.485 ;
        RECT 25.070 119.950 25.240 120.120 ;
        RECT 25.070 119.540 25.240 119.710 ;
        RECT 25.860 120.315 26.030 120.485 ;
        RECT 25.860 119.950 26.030 120.120 ;
        RECT 25.860 119.540 26.030 119.710 ;
        RECT 26.650 120.315 26.820 120.485 ;
        RECT 26.650 119.950 26.820 120.120 ;
        RECT 26.650 119.540 26.820 119.710 ;
        RECT 27.440 120.315 27.610 120.485 ;
        RECT 27.440 119.950 27.610 120.120 ;
        RECT 27.440 119.540 27.610 119.710 ;
        RECT 28.230 120.315 28.400 120.485 ;
        RECT 28.230 119.950 28.400 120.120 ;
        RECT 28.230 119.540 28.400 119.710 ;
        RECT 29.020 120.315 29.190 120.485 ;
        RECT 29.020 119.950 29.190 120.120 ;
        RECT 29.020 119.540 29.190 119.710 ;
        RECT 29.810 120.315 29.980 120.485 ;
        RECT 29.810 119.950 29.980 120.120 ;
        RECT 29.810 119.540 29.980 119.710 ;
        RECT 33.305 120.315 33.475 120.485 ;
        RECT 33.305 119.950 33.475 120.120 ;
        RECT 33.305 119.540 33.475 119.710 ;
        RECT 34.095 120.315 34.265 120.485 ;
        RECT 34.095 119.950 34.265 120.120 ;
        RECT 34.095 119.540 34.265 119.710 ;
        RECT 34.885 120.315 35.055 120.485 ;
        RECT 34.885 119.950 35.055 120.120 ;
        RECT 34.885 119.540 35.055 119.710 ;
        RECT 35.675 120.315 35.845 120.485 ;
        RECT 35.675 119.950 35.845 120.120 ;
        RECT 35.675 119.540 35.845 119.710 ;
        RECT 36.465 120.315 36.635 120.485 ;
        RECT 36.465 119.950 36.635 120.120 ;
        RECT 36.465 119.540 36.635 119.710 ;
        RECT 37.255 120.315 37.425 120.485 ;
        RECT 37.255 119.950 37.425 120.120 ;
        RECT 37.255 119.540 37.425 119.710 ;
        RECT 38.045 120.315 38.215 120.485 ;
        RECT 38.045 119.950 38.215 120.120 ;
        RECT 38.045 119.540 38.215 119.710 ;
        RECT 38.835 120.315 39.005 120.485 ;
        RECT 38.835 119.950 39.005 120.120 ;
        RECT 38.835 119.540 39.005 119.710 ;
        RECT 39.625 120.315 39.795 120.485 ;
        RECT 39.625 119.950 39.795 120.120 ;
        RECT 39.625 119.540 39.795 119.710 ;
        RECT 40.415 120.315 40.585 120.485 ;
        RECT 40.415 119.950 40.585 120.120 ;
        RECT 40.415 119.540 40.585 119.710 ;
        RECT 41.205 120.315 41.375 120.485 ;
        RECT 41.205 119.950 41.375 120.120 ;
        RECT 41.205 119.540 41.375 119.710 ;
        RECT 41.995 120.315 42.165 120.485 ;
        RECT 41.995 119.950 42.165 120.120 ;
        RECT 41.995 119.540 42.165 119.710 ;
        RECT 42.785 120.315 42.955 120.485 ;
        RECT 42.785 119.950 42.955 120.120 ;
        RECT 42.785 119.540 42.955 119.710 ;
        RECT 43.575 120.315 43.745 120.485 ;
        RECT 43.575 119.950 43.745 120.120 ;
        RECT 43.575 119.540 43.745 119.710 ;
        RECT 44.365 120.315 44.535 120.485 ;
        RECT 44.365 119.950 44.535 120.120 ;
        RECT 44.365 119.540 44.535 119.710 ;
        RECT 45.155 120.315 45.325 120.485 ;
        RECT 45.155 119.950 45.325 120.120 ;
        RECT 45.155 119.540 45.325 119.710 ;
        RECT 45.945 120.315 46.115 120.485 ;
        RECT 45.945 119.950 46.115 120.120 ;
        RECT 45.945 119.540 46.115 119.710 ;
        RECT 46.735 120.315 46.905 120.485 ;
        RECT 46.735 119.950 46.905 120.120 ;
        RECT 46.735 119.540 46.905 119.710 ;
        RECT 47.525 120.315 47.695 120.485 ;
        RECT 47.525 119.950 47.695 120.120 ;
        RECT 47.525 119.540 47.695 119.710 ;
        RECT 48.315 120.315 48.485 120.485 ;
        RECT 48.315 119.950 48.485 120.120 ;
        RECT 48.315 119.540 48.485 119.710 ;
        RECT 49.105 120.315 49.275 120.485 ;
        RECT 49.105 119.950 49.275 120.120 ;
        RECT 49.105 119.540 49.275 119.710 ;
        RECT 49.895 120.315 50.065 120.485 ;
        RECT 49.895 119.950 50.065 120.120 ;
        RECT 49.895 119.540 50.065 119.710 ;
        RECT 55.005 118.350 55.175 118.520 ;
        RECT 55.485 118.350 55.655 118.520 ;
        RECT 55.955 118.350 56.125 118.520 ;
        RECT 56.435 118.350 56.605 118.520 ;
        RECT 56.975 118.350 57.145 118.520 ;
        RECT 57.455 118.350 57.625 118.520 ;
        RECT 57.930 118.350 58.100 118.520 ;
        RECT 58.410 118.350 58.580 118.520 ;
        RECT 58.970 118.350 59.140 118.520 ;
        RECT 55.005 117.990 55.175 118.160 ;
        RECT 55.485 117.990 55.655 118.160 ;
        RECT 55.955 117.990 56.125 118.160 ;
        RECT 56.435 117.990 56.605 118.160 ;
        RECT 56.975 117.990 57.145 118.160 ;
        RECT 57.455 117.990 57.625 118.160 ;
        RECT 57.930 117.990 58.100 118.160 ;
        RECT 58.410 117.990 58.580 118.160 ;
        RECT 58.970 117.990 59.140 118.160 ;
        RECT 55.005 117.630 55.175 117.800 ;
        RECT 55.485 117.630 55.655 117.800 ;
        RECT 55.955 117.630 56.125 117.800 ;
        RECT 56.435 117.630 56.605 117.800 ;
        RECT 56.975 117.630 57.145 117.800 ;
        RECT 57.455 117.630 57.625 117.800 ;
        RECT 57.930 117.630 58.100 117.800 ;
        RECT 58.410 117.630 58.580 117.800 ;
        RECT 58.970 117.630 59.140 117.800 ;
        RECT 62.935 118.350 63.105 118.520 ;
        RECT 63.415 118.350 63.585 118.520 ;
        RECT 63.885 118.350 64.055 118.520 ;
        RECT 64.365 118.350 64.535 118.520 ;
        RECT 64.905 118.350 65.075 118.520 ;
        RECT 65.385 118.350 65.555 118.520 ;
        RECT 65.860 118.350 66.030 118.520 ;
        RECT 66.340 118.350 66.510 118.520 ;
        RECT 66.900 118.350 67.070 118.520 ;
        RECT 67.380 118.350 67.550 118.520 ;
        RECT 67.855 118.350 68.025 118.520 ;
        RECT 68.335 118.350 68.505 118.520 ;
        RECT 68.875 118.350 69.045 118.520 ;
        RECT 69.355 118.350 69.525 118.520 ;
        RECT 62.935 117.990 63.105 118.160 ;
        RECT 63.415 117.990 63.585 118.160 ;
        RECT 63.885 117.990 64.055 118.160 ;
        RECT 64.365 117.990 64.535 118.160 ;
        RECT 64.905 117.990 65.075 118.160 ;
        RECT 65.385 117.990 65.555 118.160 ;
        RECT 65.860 117.990 66.030 118.160 ;
        RECT 66.340 117.990 66.510 118.160 ;
        RECT 66.900 117.990 67.070 118.160 ;
        RECT 67.380 117.990 67.550 118.160 ;
        RECT 67.855 117.990 68.025 118.160 ;
        RECT 68.335 117.990 68.505 118.160 ;
        RECT 68.875 117.990 69.045 118.160 ;
        RECT 69.355 117.990 69.525 118.160 ;
        RECT 62.935 117.630 63.105 117.800 ;
        RECT 63.415 117.630 63.585 117.800 ;
        RECT 63.885 117.630 64.055 117.800 ;
        RECT 64.365 117.630 64.535 117.800 ;
        RECT 64.905 117.630 65.075 117.800 ;
        RECT 65.385 117.630 65.555 117.800 ;
        RECT 65.860 117.630 66.030 117.800 ;
        RECT 66.340 117.630 66.510 117.800 ;
        RECT 66.900 117.630 67.070 117.800 ;
        RECT 67.380 117.630 67.550 117.800 ;
        RECT 67.855 117.630 68.025 117.800 ;
        RECT 68.335 117.630 68.505 117.800 ;
        RECT 68.875 117.630 69.045 117.800 ;
        RECT 69.355 117.630 69.525 117.800 ;
        RECT 55.005 111.620 55.175 111.790 ;
        RECT 55.485 111.620 55.655 111.790 ;
        RECT 55.955 111.620 56.125 111.790 ;
        RECT 56.435 111.620 56.605 111.790 ;
        RECT 56.975 111.620 57.145 111.790 ;
        RECT 57.455 111.620 57.625 111.790 ;
        RECT 57.930 111.620 58.100 111.790 ;
        RECT 58.410 111.620 58.580 111.790 ;
        RECT 58.970 111.620 59.140 111.790 ;
        RECT 55.005 111.260 55.175 111.430 ;
        RECT 55.485 111.260 55.655 111.430 ;
        RECT 55.955 111.260 56.125 111.430 ;
        RECT 56.435 111.260 56.605 111.430 ;
        RECT 56.975 111.260 57.145 111.430 ;
        RECT 57.455 111.260 57.625 111.430 ;
        RECT 57.930 111.260 58.100 111.430 ;
        RECT 58.410 111.260 58.580 111.430 ;
        RECT 58.970 111.260 59.140 111.430 ;
        RECT 55.005 110.900 55.175 111.070 ;
        RECT 55.485 110.900 55.655 111.070 ;
        RECT 55.955 110.900 56.125 111.070 ;
        RECT 56.435 110.900 56.605 111.070 ;
        RECT 56.975 110.900 57.145 111.070 ;
        RECT 57.455 110.900 57.625 111.070 ;
        RECT 57.930 110.900 58.100 111.070 ;
        RECT 58.410 110.900 58.580 111.070 ;
        RECT 58.970 110.900 59.140 111.070 ;
        RECT 62.935 111.620 63.105 111.790 ;
        RECT 63.415 111.620 63.585 111.790 ;
        RECT 63.885 111.620 64.055 111.790 ;
        RECT 64.365 111.620 64.535 111.790 ;
        RECT 64.905 111.620 65.075 111.790 ;
        RECT 65.385 111.620 65.555 111.790 ;
        RECT 65.860 111.620 66.030 111.790 ;
        RECT 66.340 111.620 66.510 111.790 ;
        RECT 66.900 111.620 67.070 111.790 ;
        RECT 67.380 111.620 67.550 111.790 ;
        RECT 67.855 111.620 68.025 111.790 ;
        RECT 68.335 111.620 68.505 111.790 ;
        RECT 68.875 111.620 69.045 111.790 ;
        RECT 69.355 111.620 69.525 111.790 ;
        RECT 62.935 111.260 63.105 111.430 ;
        RECT 63.415 111.260 63.585 111.430 ;
        RECT 63.885 111.260 64.055 111.430 ;
        RECT 64.365 111.260 64.535 111.430 ;
        RECT 64.905 111.260 65.075 111.430 ;
        RECT 65.385 111.260 65.555 111.430 ;
        RECT 65.860 111.260 66.030 111.430 ;
        RECT 66.340 111.260 66.510 111.430 ;
        RECT 66.900 111.260 67.070 111.430 ;
        RECT 67.380 111.260 67.550 111.430 ;
        RECT 67.855 111.260 68.025 111.430 ;
        RECT 68.335 111.260 68.505 111.430 ;
        RECT 68.875 111.260 69.045 111.430 ;
        RECT 69.355 111.260 69.525 111.430 ;
        RECT 62.935 110.900 63.105 111.070 ;
        RECT 63.415 110.900 63.585 111.070 ;
        RECT 63.885 110.900 64.055 111.070 ;
        RECT 64.365 110.900 64.535 111.070 ;
        RECT 64.905 110.900 65.075 111.070 ;
        RECT 65.385 110.900 65.555 111.070 ;
        RECT 65.860 110.900 66.030 111.070 ;
        RECT 66.340 110.900 66.510 111.070 ;
        RECT 66.900 110.900 67.070 111.070 ;
        RECT 67.380 110.900 67.550 111.070 ;
        RECT 67.855 110.900 68.025 111.070 ;
        RECT 68.335 110.900 68.505 111.070 ;
        RECT 68.875 110.900 69.045 111.070 ;
        RECT 69.355 110.900 69.525 111.070 ;
        RECT 16.460 108.510 16.630 108.680 ;
        RECT 16.460 108.060 16.630 108.230 ;
        RECT 16.460 107.670 16.630 107.840 ;
        RECT 17.250 108.510 17.420 108.680 ;
        RECT 17.250 108.060 17.420 108.230 ;
        RECT 17.250 107.670 17.420 107.840 ;
        RECT 18.040 108.510 18.210 108.680 ;
        RECT 18.040 108.060 18.210 108.230 ;
        RECT 18.040 107.670 18.210 107.840 ;
        RECT 18.830 108.510 19.000 108.680 ;
        RECT 18.830 108.060 19.000 108.230 ;
        RECT 18.830 107.670 19.000 107.840 ;
        RECT 19.620 108.510 19.790 108.680 ;
        RECT 19.620 108.060 19.790 108.230 ;
        RECT 19.620 107.670 19.790 107.840 ;
        RECT 20.410 108.510 20.580 108.680 ;
        RECT 20.410 108.060 20.580 108.230 ;
        RECT 20.410 107.670 20.580 107.840 ;
        RECT 23.490 108.510 23.660 108.680 ;
        RECT 23.490 108.060 23.660 108.230 ;
        RECT 23.490 107.670 23.660 107.840 ;
        RECT 24.280 108.510 24.450 108.680 ;
        RECT 24.280 108.060 24.450 108.230 ;
        RECT 24.280 107.670 24.450 107.840 ;
        RECT 25.070 108.510 25.240 108.680 ;
        RECT 25.070 108.060 25.240 108.230 ;
        RECT 25.070 107.670 25.240 107.840 ;
        RECT 25.860 108.510 26.030 108.680 ;
        RECT 25.860 108.060 26.030 108.230 ;
        RECT 25.860 107.670 26.030 107.840 ;
        RECT 26.650 108.510 26.820 108.680 ;
        RECT 26.650 108.060 26.820 108.230 ;
        RECT 26.650 107.670 26.820 107.840 ;
        RECT 27.440 108.510 27.610 108.680 ;
        RECT 27.440 108.060 27.610 108.230 ;
        RECT 27.440 107.670 27.610 107.840 ;
        RECT 28.230 108.510 28.400 108.680 ;
        RECT 28.230 108.060 28.400 108.230 ;
        RECT 28.230 107.670 28.400 107.840 ;
        RECT 29.020 108.510 29.190 108.680 ;
        RECT 29.020 108.060 29.190 108.230 ;
        RECT 29.020 107.670 29.190 107.840 ;
        RECT 29.810 108.510 29.980 108.680 ;
        RECT 29.810 108.060 29.980 108.230 ;
        RECT 29.810 107.670 29.980 107.840 ;
        RECT 33.305 108.510 33.475 108.680 ;
        RECT 33.305 108.060 33.475 108.230 ;
        RECT 33.305 107.670 33.475 107.840 ;
        RECT 34.095 108.510 34.265 108.680 ;
        RECT 34.095 108.060 34.265 108.230 ;
        RECT 34.095 107.670 34.265 107.840 ;
        RECT 34.885 108.510 35.055 108.680 ;
        RECT 34.885 108.060 35.055 108.230 ;
        RECT 34.885 107.670 35.055 107.840 ;
        RECT 35.675 108.510 35.845 108.680 ;
        RECT 35.675 108.060 35.845 108.230 ;
        RECT 35.675 107.670 35.845 107.840 ;
        RECT 36.465 108.510 36.635 108.680 ;
        RECT 36.465 108.060 36.635 108.230 ;
        RECT 36.465 107.670 36.635 107.840 ;
        RECT 37.255 108.510 37.425 108.680 ;
        RECT 37.255 108.060 37.425 108.230 ;
        RECT 37.255 107.670 37.425 107.840 ;
        RECT 38.045 108.510 38.215 108.680 ;
        RECT 38.045 108.060 38.215 108.230 ;
        RECT 38.045 107.670 38.215 107.840 ;
        RECT 38.835 108.510 39.005 108.680 ;
        RECT 38.835 108.060 39.005 108.230 ;
        RECT 38.835 107.670 39.005 107.840 ;
        RECT 39.625 108.510 39.795 108.680 ;
        RECT 39.625 108.060 39.795 108.230 ;
        RECT 39.625 107.670 39.795 107.840 ;
        RECT 40.415 108.510 40.585 108.680 ;
        RECT 40.415 108.060 40.585 108.230 ;
        RECT 40.415 107.670 40.585 107.840 ;
        RECT 41.205 108.510 41.375 108.680 ;
        RECT 41.205 108.060 41.375 108.230 ;
        RECT 41.205 107.670 41.375 107.840 ;
        RECT 41.995 108.510 42.165 108.680 ;
        RECT 41.995 108.060 42.165 108.230 ;
        RECT 41.995 107.670 42.165 107.840 ;
        RECT 42.785 108.510 42.955 108.680 ;
        RECT 42.785 108.060 42.955 108.230 ;
        RECT 42.785 107.670 42.955 107.840 ;
        RECT 43.575 108.510 43.745 108.680 ;
        RECT 43.575 108.060 43.745 108.230 ;
        RECT 43.575 107.670 43.745 107.840 ;
        RECT 44.365 108.510 44.535 108.680 ;
        RECT 44.365 108.060 44.535 108.230 ;
        RECT 44.365 107.670 44.535 107.840 ;
        RECT 45.155 108.510 45.325 108.680 ;
        RECT 45.155 108.060 45.325 108.230 ;
        RECT 45.155 107.670 45.325 107.840 ;
        RECT 45.945 108.510 46.115 108.680 ;
        RECT 45.945 108.060 46.115 108.230 ;
        RECT 45.945 107.670 46.115 107.840 ;
        RECT 46.735 108.510 46.905 108.680 ;
        RECT 46.735 108.060 46.905 108.230 ;
        RECT 46.735 107.670 46.905 107.840 ;
        RECT 47.525 108.510 47.695 108.680 ;
        RECT 47.525 108.060 47.695 108.230 ;
        RECT 47.525 107.670 47.695 107.840 ;
        RECT 48.315 108.510 48.485 108.680 ;
        RECT 48.315 108.060 48.485 108.230 ;
        RECT 48.315 107.670 48.485 107.840 ;
        RECT 49.105 108.510 49.275 108.680 ;
        RECT 49.105 108.060 49.275 108.230 ;
        RECT 49.105 107.670 49.275 107.840 ;
        RECT 49.895 108.510 50.065 108.680 ;
        RECT 49.895 108.060 50.065 108.230 ;
        RECT 49.895 107.670 50.065 107.840 ;
        RECT 20.160 104.315 20.330 104.485 ;
        RECT 15.720 103.575 15.890 103.745 ;
        RECT 16.080 103.575 16.250 103.745 ;
        RECT 18.445 103.700 18.615 103.870 ;
        RECT 18.805 103.700 18.975 103.870 ;
        RECT 21.720 104.315 21.890 104.485 ;
        RECT 20.770 103.575 20.940 103.745 ;
        RECT 21.130 103.575 21.300 103.745 ;
        RECT 23.280 104.315 23.450 104.485 ;
        RECT 22.320 103.575 22.490 103.745 ;
        RECT 22.680 103.575 22.850 103.745 ;
        RECT 24.840 104.315 25.010 104.485 ;
        RECT 23.880 103.575 24.050 103.745 ;
        RECT 24.240 103.575 24.410 103.745 ;
        RECT 26.400 104.315 26.570 104.485 ;
        RECT 25.440 103.575 25.610 103.745 ;
        RECT 25.800 103.575 25.970 103.745 ;
        RECT 27.960 104.315 28.130 104.485 ;
        RECT 27.000 103.575 27.170 103.745 ;
        RECT 27.360 103.575 27.530 103.745 ;
        RECT 29.520 104.315 29.690 104.485 ;
        RECT 28.560 103.575 28.730 103.745 ;
        RECT 28.920 103.575 29.090 103.745 ;
        RECT 31.080 104.315 31.250 104.485 ;
        RECT 30.120 103.575 30.290 103.745 ;
        RECT 30.480 103.575 30.650 103.745 ;
        RECT 37.440 104.315 37.610 104.485 ;
        RECT 32.820 103.575 32.990 103.745 ;
        RECT 33.180 103.575 33.350 103.745 ;
        RECT 35.725 103.700 35.895 103.870 ;
        RECT 36.085 103.700 36.255 103.870 ;
        RECT 39.000 104.315 39.170 104.485 ;
        RECT 38.050 103.575 38.220 103.745 ;
        RECT 38.410 103.575 38.580 103.745 ;
        RECT 40.560 104.315 40.730 104.485 ;
        RECT 39.600 103.575 39.770 103.745 ;
        RECT 39.960 103.575 40.130 103.745 ;
        RECT 42.120 104.315 42.290 104.485 ;
        RECT 41.160 103.575 41.330 103.745 ;
        RECT 41.520 103.575 41.690 103.745 ;
        RECT 43.680 104.315 43.850 104.485 ;
        RECT 42.720 103.575 42.890 103.745 ;
        RECT 43.080 103.575 43.250 103.745 ;
        RECT 45.240 104.315 45.410 104.485 ;
        RECT 44.280 103.575 44.450 103.745 ;
        RECT 44.640 103.575 44.810 103.745 ;
        RECT 46.800 104.315 46.970 104.485 ;
        RECT 45.840 103.575 46.010 103.745 ;
        RECT 46.200 103.575 46.370 103.745 ;
        RECT 48.360 104.315 48.530 104.485 ;
        RECT 47.400 103.575 47.570 103.745 ;
        RECT 47.760 103.575 47.930 103.745 ;
        RECT 54.720 104.315 54.890 104.485 ;
        RECT 50.250 103.575 50.420 103.745 ;
        RECT 50.610 103.575 50.780 103.745 ;
        RECT 52.995 103.700 53.165 103.870 ;
        RECT 53.355 103.700 53.525 103.870 ;
        RECT 56.280 104.315 56.450 104.485 ;
        RECT 55.330 103.575 55.500 103.745 ;
        RECT 55.690 103.575 55.860 103.745 ;
        RECT 57.840 104.315 58.010 104.485 ;
        RECT 56.880 103.575 57.050 103.745 ;
        RECT 57.240 103.575 57.410 103.745 ;
        RECT 59.400 104.315 59.570 104.485 ;
        RECT 58.440 103.575 58.610 103.745 ;
        RECT 58.800 103.575 58.970 103.745 ;
        RECT 60.960 104.315 61.130 104.485 ;
        RECT 60.000 103.575 60.170 103.745 ;
        RECT 60.360 103.575 60.530 103.745 ;
        RECT 62.520 104.315 62.690 104.485 ;
        RECT 61.560 103.575 61.730 103.745 ;
        RECT 61.920 103.575 62.090 103.745 ;
        RECT 64.080 104.315 64.250 104.485 ;
        RECT 63.120 103.575 63.290 103.745 ;
        RECT 63.480 103.575 63.650 103.745 ;
        RECT 65.640 104.315 65.810 104.485 ;
        RECT 64.680 103.575 64.850 103.745 ;
        RECT 65.040 103.575 65.210 103.745 ;
        RECT 15.720 100.245 15.890 100.415 ;
        RECT 16.080 100.245 16.250 100.415 ;
        RECT 18.445 100.080 18.615 100.250 ;
        RECT 18.805 100.080 18.975 100.250 ;
        RECT 20.770 100.245 20.940 100.415 ;
        RECT 21.130 100.245 21.300 100.415 ;
        RECT 20.160 99.505 20.330 99.675 ;
        RECT 22.320 100.245 22.490 100.415 ;
        RECT 22.680 100.245 22.850 100.415 ;
        RECT 21.720 99.505 21.890 99.675 ;
        RECT 23.880 100.245 24.050 100.415 ;
        RECT 24.240 100.245 24.410 100.415 ;
        RECT 23.280 99.505 23.450 99.675 ;
        RECT 25.440 100.245 25.610 100.415 ;
        RECT 25.800 100.245 25.970 100.415 ;
        RECT 24.840 99.505 25.010 99.675 ;
        RECT 27.000 100.245 27.170 100.415 ;
        RECT 27.360 100.245 27.530 100.415 ;
        RECT 26.400 99.505 26.570 99.675 ;
        RECT 28.560 100.245 28.730 100.415 ;
        RECT 28.920 100.245 29.090 100.415 ;
        RECT 27.960 99.505 28.130 99.675 ;
        RECT 30.120 100.245 30.290 100.415 ;
        RECT 30.480 100.245 30.650 100.415 ;
        RECT 29.520 99.505 29.690 99.675 ;
        RECT 32.975 100.245 33.145 100.415 ;
        RECT 33.335 100.245 33.505 100.415 ;
        RECT 35.725 100.085 35.895 100.255 ;
        RECT 36.085 100.085 36.255 100.255 ;
        RECT 31.080 99.505 31.250 99.675 ;
        RECT 38.050 100.245 38.220 100.415 ;
        RECT 38.410 100.245 38.580 100.415 ;
        RECT 37.440 99.505 37.610 99.675 ;
        RECT 39.600 100.245 39.770 100.415 ;
        RECT 39.960 100.245 40.130 100.415 ;
        RECT 39.000 99.505 39.170 99.675 ;
        RECT 41.160 100.245 41.330 100.415 ;
        RECT 41.520 100.245 41.690 100.415 ;
        RECT 40.560 99.505 40.730 99.675 ;
        RECT 42.720 100.245 42.890 100.415 ;
        RECT 43.080 100.245 43.250 100.415 ;
        RECT 42.120 99.505 42.290 99.675 ;
        RECT 44.280 100.245 44.450 100.415 ;
        RECT 44.640 100.245 44.810 100.415 ;
        RECT 43.680 99.505 43.850 99.675 ;
        RECT 45.840 100.245 46.010 100.415 ;
        RECT 46.200 100.245 46.370 100.415 ;
        RECT 45.240 99.505 45.410 99.675 ;
        RECT 47.400 100.245 47.570 100.415 ;
        RECT 47.760 100.245 47.930 100.415 ;
        RECT 46.800 99.505 46.970 99.675 ;
        RECT 50.265 100.245 50.435 100.415 ;
        RECT 50.625 100.245 50.795 100.415 ;
        RECT 52.995 100.100 53.165 100.270 ;
        RECT 53.355 100.100 53.525 100.270 ;
        RECT 48.360 99.505 48.530 99.675 ;
        RECT 55.330 100.245 55.500 100.415 ;
        RECT 55.690 100.245 55.860 100.415 ;
        RECT 54.720 99.505 54.890 99.675 ;
        RECT 56.880 100.245 57.050 100.415 ;
        RECT 57.240 100.245 57.410 100.415 ;
        RECT 56.280 99.505 56.450 99.675 ;
        RECT 58.440 100.245 58.610 100.415 ;
        RECT 58.800 100.245 58.970 100.415 ;
        RECT 57.840 99.505 58.010 99.675 ;
        RECT 60.000 100.245 60.170 100.415 ;
        RECT 60.360 100.245 60.530 100.415 ;
        RECT 59.400 99.505 59.570 99.675 ;
        RECT 61.560 100.245 61.730 100.415 ;
        RECT 61.920 100.245 62.090 100.415 ;
        RECT 60.960 99.505 61.130 99.675 ;
        RECT 63.120 100.245 63.290 100.415 ;
        RECT 63.480 100.245 63.650 100.415 ;
        RECT 62.520 99.505 62.690 99.675 ;
        RECT 64.680 100.245 64.850 100.415 ;
        RECT 65.040 100.245 65.210 100.415 ;
        RECT 64.080 99.505 64.250 99.675 ;
        RECT 65.640 99.505 65.810 99.675 ;
        RECT 16.845 95.885 17.015 96.055 ;
        RECT 17.205 95.885 17.375 96.055 ;
        RECT 19.575 95.885 19.745 96.055 ;
        RECT 19.935 95.885 20.105 96.055 ;
        RECT 22.605 95.885 22.775 96.055 ;
        RECT 22.965 95.885 23.135 96.055 ;
        RECT 25.335 95.885 25.505 96.055 ;
        RECT 25.695 95.885 25.865 96.055 ;
        RECT 28.365 95.885 28.535 96.055 ;
        RECT 28.725 95.885 28.895 96.055 ;
        RECT 31.095 95.885 31.265 96.055 ;
        RECT 31.455 95.885 31.625 96.055 ;
        RECT 34.125 95.885 34.295 96.055 ;
        RECT 34.485 95.885 34.655 96.055 ;
        RECT 36.855 95.885 37.025 96.055 ;
        RECT 37.215 95.885 37.385 96.055 ;
        RECT 39.885 95.885 40.055 96.055 ;
        RECT 40.245 95.885 40.415 96.055 ;
        RECT 42.615 95.885 42.785 96.055 ;
        RECT 42.975 95.885 43.145 96.055 ;
        RECT 45.645 95.885 45.815 96.055 ;
        RECT 46.005 95.885 46.175 96.055 ;
        RECT 48.375 95.885 48.545 96.055 ;
        RECT 48.735 95.885 48.905 96.055 ;
        RECT 16.845 95.095 17.015 95.265 ;
        RECT 17.205 95.095 17.375 95.265 ;
        RECT 19.575 95.095 19.745 95.265 ;
        RECT 19.935 95.095 20.105 95.265 ;
        RECT 22.605 95.095 22.775 95.265 ;
        RECT 22.965 95.095 23.135 95.265 ;
        RECT 25.335 95.095 25.505 95.265 ;
        RECT 25.695 95.095 25.865 95.265 ;
        RECT 28.365 95.095 28.535 95.265 ;
        RECT 28.725 95.095 28.895 95.265 ;
        RECT 31.095 95.095 31.265 95.265 ;
        RECT 31.455 95.095 31.625 95.265 ;
        RECT 34.125 95.095 34.295 95.265 ;
        RECT 34.485 95.095 34.655 95.265 ;
        RECT 36.855 95.095 37.025 95.265 ;
        RECT 37.215 95.095 37.385 95.265 ;
        RECT 39.885 95.095 40.055 95.265 ;
        RECT 40.245 95.095 40.415 95.265 ;
        RECT 42.615 95.095 42.785 95.265 ;
        RECT 42.975 95.095 43.145 95.265 ;
        RECT 45.645 95.095 45.815 95.265 ;
        RECT 46.005 95.095 46.175 95.265 ;
        RECT 48.375 95.095 48.545 95.265 ;
        RECT 48.735 95.095 48.905 95.265 ;
        RECT 18.330 94.700 18.500 94.870 ;
        RECT 18.690 94.700 18.860 94.870 ;
        RECT 24.090 94.700 24.260 94.870 ;
        RECT 24.450 94.700 24.620 94.870 ;
        RECT 29.850 94.700 30.020 94.870 ;
        RECT 30.210 94.700 30.380 94.870 ;
        RECT 35.610 94.700 35.780 94.870 ;
        RECT 35.970 94.700 36.140 94.870 ;
        RECT 41.370 94.700 41.540 94.870 ;
        RECT 41.730 94.700 41.900 94.870 ;
        RECT 47.130 94.700 47.300 94.870 ;
        RECT 47.490 94.700 47.660 94.870 ;
        RECT 52.930 94.275 53.100 94.445 ;
        RECT 53.410 94.275 53.580 94.445 ;
        RECT 53.880 94.275 54.050 94.445 ;
        RECT 54.360 94.275 54.530 94.445 ;
        RECT 54.900 94.275 55.070 94.445 ;
        RECT 55.380 94.275 55.550 94.445 ;
        RECT 55.855 94.275 56.025 94.445 ;
        RECT 56.335 94.275 56.505 94.445 ;
        RECT 56.895 94.275 57.065 94.445 ;
        RECT 57.375 94.275 57.545 94.445 ;
        RECT 57.850 94.275 58.020 94.445 ;
        RECT 58.330 94.275 58.500 94.445 ;
        RECT 58.870 94.275 59.040 94.445 ;
        RECT 59.350 94.275 59.520 94.445 ;
        RECT 59.825 94.275 59.995 94.445 ;
        RECT 60.305 94.275 60.475 94.445 ;
        RECT 60.895 94.275 61.065 94.445 ;
        RECT 61.375 94.275 61.545 94.445 ;
        RECT 61.850 94.275 62.020 94.445 ;
        RECT 62.330 94.275 62.500 94.445 ;
        RECT 62.870 94.275 63.040 94.445 ;
        RECT 63.350 94.275 63.520 94.445 ;
        RECT 63.825 94.275 63.995 94.445 ;
        RECT 64.305 94.275 64.475 94.445 ;
        RECT 64.865 94.275 65.035 94.445 ;
        RECT 65.345 94.275 65.515 94.445 ;
        RECT 65.820 94.275 65.990 94.445 ;
        RECT 66.300 94.275 66.470 94.445 ;
        RECT 66.840 94.275 67.010 94.445 ;
        RECT 67.320 94.275 67.490 94.445 ;
        RECT 67.795 94.275 67.965 94.445 ;
        RECT 68.275 94.275 68.445 94.445 ;
        RECT 52.930 93.915 53.100 94.085 ;
        RECT 53.410 93.915 53.580 94.085 ;
        RECT 53.880 93.915 54.050 94.085 ;
        RECT 54.360 93.915 54.530 94.085 ;
        RECT 54.900 93.915 55.070 94.085 ;
        RECT 55.380 93.915 55.550 94.085 ;
        RECT 55.855 93.915 56.025 94.085 ;
        RECT 56.335 93.915 56.505 94.085 ;
        RECT 56.895 93.915 57.065 94.085 ;
        RECT 57.375 93.915 57.545 94.085 ;
        RECT 57.850 93.915 58.020 94.085 ;
        RECT 58.330 93.915 58.500 94.085 ;
        RECT 58.870 93.915 59.040 94.085 ;
        RECT 59.350 93.915 59.520 94.085 ;
        RECT 59.825 93.915 59.995 94.085 ;
        RECT 60.305 93.915 60.475 94.085 ;
        RECT 60.895 93.915 61.065 94.085 ;
        RECT 61.375 93.915 61.545 94.085 ;
        RECT 61.850 93.915 62.020 94.085 ;
        RECT 62.330 93.915 62.500 94.085 ;
        RECT 62.870 93.915 63.040 94.085 ;
        RECT 63.350 93.915 63.520 94.085 ;
        RECT 63.825 93.915 63.995 94.085 ;
        RECT 64.305 93.915 64.475 94.085 ;
        RECT 64.865 93.915 65.035 94.085 ;
        RECT 65.345 93.915 65.515 94.085 ;
        RECT 65.820 93.915 65.990 94.085 ;
        RECT 66.300 93.915 66.470 94.085 ;
        RECT 66.840 93.915 67.010 94.085 ;
        RECT 67.320 93.915 67.490 94.085 ;
        RECT 67.795 93.915 67.965 94.085 ;
        RECT 68.275 93.915 68.445 94.085 ;
        RECT 16.765 93.480 16.935 93.650 ;
        RECT 17.125 93.480 17.295 93.650 ;
        RECT 19.560 93.480 19.730 93.650 ;
        RECT 19.920 93.480 20.090 93.650 ;
        RECT 22.525 93.480 22.695 93.650 ;
        RECT 22.885 93.480 23.055 93.650 ;
        RECT 25.320 93.480 25.490 93.650 ;
        RECT 25.680 93.480 25.850 93.650 ;
        RECT 28.285 93.480 28.455 93.650 ;
        RECT 28.645 93.480 28.815 93.650 ;
        RECT 31.080 93.480 31.250 93.650 ;
        RECT 31.440 93.480 31.610 93.650 ;
        RECT 34.045 93.480 34.215 93.650 ;
        RECT 34.405 93.480 34.575 93.650 ;
        RECT 36.840 93.480 37.010 93.650 ;
        RECT 37.200 93.480 37.370 93.650 ;
        RECT 39.805 93.480 39.975 93.650 ;
        RECT 40.165 93.480 40.335 93.650 ;
        RECT 42.600 93.480 42.770 93.650 ;
        RECT 42.960 93.480 43.130 93.650 ;
        RECT 45.565 93.480 45.735 93.650 ;
        RECT 45.925 93.480 46.095 93.650 ;
        RECT 48.360 93.480 48.530 93.650 ;
        RECT 48.720 93.480 48.890 93.650 ;
        RECT 52.930 93.555 53.100 93.725 ;
        RECT 53.410 93.555 53.580 93.725 ;
        RECT 53.880 93.555 54.050 93.725 ;
        RECT 54.360 93.555 54.530 93.725 ;
        RECT 54.900 93.555 55.070 93.725 ;
        RECT 55.380 93.555 55.550 93.725 ;
        RECT 55.855 93.555 56.025 93.725 ;
        RECT 56.335 93.555 56.505 93.725 ;
        RECT 56.895 93.555 57.065 93.725 ;
        RECT 57.375 93.555 57.545 93.725 ;
        RECT 57.850 93.555 58.020 93.725 ;
        RECT 58.330 93.555 58.500 93.725 ;
        RECT 58.870 93.555 59.040 93.725 ;
        RECT 59.350 93.555 59.520 93.725 ;
        RECT 59.825 93.555 59.995 93.725 ;
        RECT 60.305 93.555 60.475 93.725 ;
        RECT 60.895 93.555 61.065 93.725 ;
        RECT 61.375 93.555 61.545 93.725 ;
        RECT 61.850 93.555 62.020 93.725 ;
        RECT 62.330 93.555 62.500 93.725 ;
        RECT 62.870 93.555 63.040 93.725 ;
        RECT 63.350 93.555 63.520 93.725 ;
        RECT 63.825 93.555 63.995 93.725 ;
        RECT 64.305 93.555 64.475 93.725 ;
        RECT 64.865 93.555 65.035 93.725 ;
        RECT 65.345 93.555 65.515 93.725 ;
        RECT 65.820 93.555 65.990 93.725 ;
        RECT 66.300 93.555 66.470 93.725 ;
        RECT 66.840 93.555 67.010 93.725 ;
        RECT 67.320 93.555 67.490 93.725 ;
        RECT 67.795 93.555 67.965 93.725 ;
        RECT 68.275 93.555 68.445 93.725 ;
        RECT 18.270 92.145 18.440 92.315 ;
        RECT 18.630 92.145 18.800 92.315 ;
        RECT 24.030 92.145 24.200 92.315 ;
        RECT 24.390 92.145 24.560 92.315 ;
        RECT 29.790 92.145 29.960 92.315 ;
        RECT 30.150 92.145 30.320 92.315 ;
        RECT 35.550 92.145 35.720 92.315 ;
        RECT 35.910 92.145 36.080 92.315 ;
        RECT 41.310 92.145 41.480 92.315 ;
        RECT 41.670 92.145 41.840 92.315 ;
        RECT 47.070 92.145 47.240 92.315 ;
        RECT 47.430 92.145 47.600 92.315 ;
        RECT 16.835 91.815 17.005 91.985 ;
        RECT 17.195 91.815 17.365 91.985 ;
        RECT 19.465 91.750 19.635 91.920 ;
        RECT 19.825 91.750 19.995 91.920 ;
        RECT 22.595 91.815 22.765 91.985 ;
        RECT 22.955 91.815 23.125 91.985 ;
        RECT 25.225 91.750 25.395 91.920 ;
        RECT 25.585 91.750 25.755 91.920 ;
        RECT 28.355 91.815 28.525 91.985 ;
        RECT 28.715 91.815 28.885 91.985 ;
        RECT 30.985 91.750 31.155 91.920 ;
        RECT 31.345 91.750 31.515 91.920 ;
        RECT 34.115 91.815 34.285 91.985 ;
        RECT 34.475 91.815 34.645 91.985 ;
        RECT 36.745 91.750 36.915 91.920 ;
        RECT 37.105 91.750 37.275 91.920 ;
        RECT 39.875 91.815 40.045 91.985 ;
        RECT 40.235 91.815 40.405 91.985 ;
        RECT 42.505 91.750 42.675 91.920 ;
        RECT 42.865 91.750 43.035 91.920 ;
        RECT 45.635 91.815 45.805 91.985 ;
        RECT 45.995 91.815 46.165 91.985 ;
        RECT 48.265 91.750 48.435 91.920 ;
        RECT 48.625 91.750 48.795 91.920 ;
        RECT 16.835 90.605 17.005 90.775 ;
        RECT 17.195 90.605 17.365 90.775 ;
        RECT 19.465 90.670 19.635 90.840 ;
        RECT 19.825 90.670 19.995 90.840 ;
        RECT 22.595 90.605 22.765 90.775 ;
        RECT 22.955 90.605 23.125 90.775 ;
        RECT 25.225 90.670 25.395 90.840 ;
        RECT 25.585 90.670 25.755 90.840 ;
        RECT 28.355 90.605 28.525 90.775 ;
        RECT 28.715 90.605 28.885 90.775 ;
        RECT 30.985 90.670 31.155 90.840 ;
        RECT 31.345 90.670 31.515 90.840 ;
        RECT 34.115 90.605 34.285 90.775 ;
        RECT 34.475 90.605 34.645 90.775 ;
        RECT 36.745 90.670 36.915 90.840 ;
        RECT 37.105 90.670 37.275 90.840 ;
        RECT 39.875 90.605 40.045 90.775 ;
        RECT 40.235 90.605 40.405 90.775 ;
        RECT 42.505 90.670 42.675 90.840 ;
        RECT 42.865 90.670 43.035 90.840 ;
        RECT 45.635 90.605 45.805 90.775 ;
        RECT 45.995 90.605 46.165 90.775 ;
        RECT 48.265 90.670 48.435 90.840 ;
        RECT 48.625 90.670 48.795 90.840 ;
        RECT 18.270 90.275 18.440 90.445 ;
        RECT 18.630 90.275 18.800 90.445 ;
        RECT 24.030 90.275 24.200 90.445 ;
        RECT 24.390 90.275 24.560 90.445 ;
        RECT 29.790 90.275 29.960 90.445 ;
        RECT 30.150 90.275 30.320 90.445 ;
        RECT 35.550 90.275 35.720 90.445 ;
        RECT 35.910 90.275 36.080 90.445 ;
        RECT 41.310 90.275 41.480 90.445 ;
        RECT 41.670 90.275 41.840 90.445 ;
        RECT 47.070 90.275 47.240 90.445 ;
        RECT 47.430 90.275 47.600 90.445 ;
        RECT 16.715 89.010 16.885 89.180 ;
        RECT 17.075 89.010 17.245 89.180 ;
        RECT 19.560 89.010 19.730 89.180 ;
        RECT 19.920 89.010 20.090 89.180 ;
        RECT 22.475 89.010 22.645 89.180 ;
        RECT 22.835 89.010 23.005 89.180 ;
        RECT 25.320 89.010 25.490 89.180 ;
        RECT 25.680 89.010 25.850 89.180 ;
        RECT 28.235 89.010 28.405 89.180 ;
        RECT 28.595 89.010 28.765 89.180 ;
        RECT 31.080 89.010 31.250 89.180 ;
        RECT 31.440 89.010 31.610 89.180 ;
        RECT 33.995 89.010 34.165 89.180 ;
        RECT 34.355 89.010 34.525 89.180 ;
        RECT 36.840 89.010 37.010 89.180 ;
        RECT 37.200 89.010 37.370 89.180 ;
        RECT 39.755 89.010 39.925 89.180 ;
        RECT 40.115 89.010 40.285 89.180 ;
        RECT 42.600 89.010 42.770 89.180 ;
        RECT 42.960 89.010 43.130 89.180 ;
        RECT 45.515 89.010 45.685 89.180 ;
        RECT 45.875 89.010 46.045 89.180 ;
        RECT 48.360 89.010 48.530 89.180 ;
        RECT 48.720 89.010 48.890 89.180 ;
        RECT 18.330 87.535 18.500 87.705 ;
        RECT 18.690 87.535 18.860 87.705 ;
        RECT 24.090 87.535 24.260 87.705 ;
        RECT 24.450 87.535 24.620 87.705 ;
        RECT 29.850 87.535 30.020 87.705 ;
        RECT 30.210 87.535 30.380 87.705 ;
        RECT 35.610 87.535 35.780 87.705 ;
        RECT 35.970 87.535 36.140 87.705 ;
        RECT 41.370 87.535 41.540 87.705 ;
        RECT 41.730 87.535 41.900 87.705 ;
        RECT 47.130 87.535 47.300 87.705 ;
        RECT 47.490 87.535 47.660 87.705 ;
        RECT 52.930 87.545 53.100 87.715 ;
        RECT 53.410 87.545 53.580 87.715 ;
        RECT 53.880 87.545 54.050 87.715 ;
        RECT 54.360 87.545 54.530 87.715 ;
        RECT 54.900 87.545 55.070 87.715 ;
        RECT 55.380 87.545 55.550 87.715 ;
        RECT 55.855 87.545 56.025 87.715 ;
        RECT 56.335 87.545 56.505 87.715 ;
        RECT 56.895 87.545 57.065 87.715 ;
        RECT 57.375 87.545 57.545 87.715 ;
        RECT 57.850 87.545 58.020 87.715 ;
        RECT 58.330 87.545 58.500 87.715 ;
        RECT 58.870 87.545 59.040 87.715 ;
        RECT 59.350 87.545 59.520 87.715 ;
        RECT 59.825 87.545 59.995 87.715 ;
        RECT 60.305 87.545 60.475 87.715 ;
        RECT 60.895 87.545 61.065 87.715 ;
        RECT 61.375 87.545 61.545 87.715 ;
        RECT 61.850 87.545 62.020 87.715 ;
        RECT 62.330 87.545 62.500 87.715 ;
        RECT 62.870 87.545 63.040 87.715 ;
        RECT 63.350 87.545 63.520 87.715 ;
        RECT 63.825 87.545 63.995 87.715 ;
        RECT 64.305 87.545 64.475 87.715 ;
        RECT 64.865 87.545 65.035 87.715 ;
        RECT 65.345 87.545 65.515 87.715 ;
        RECT 65.820 87.545 65.990 87.715 ;
        RECT 66.300 87.545 66.470 87.715 ;
        RECT 66.840 87.545 67.010 87.715 ;
        RECT 67.320 87.545 67.490 87.715 ;
        RECT 67.795 87.545 67.965 87.715 ;
        RECT 68.275 87.545 68.445 87.715 ;
        RECT 16.845 87.140 17.015 87.310 ;
        RECT 17.205 87.140 17.375 87.310 ;
        RECT 19.575 87.140 19.745 87.310 ;
        RECT 19.935 87.140 20.105 87.310 ;
        RECT 22.605 87.140 22.775 87.310 ;
        RECT 22.965 87.140 23.135 87.310 ;
        RECT 25.335 87.140 25.505 87.310 ;
        RECT 25.695 87.140 25.865 87.310 ;
        RECT 28.365 87.140 28.535 87.310 ;
        RECT 28.725 87.140 28.895 87.310 ;
        RECT 31.095 87.140 31.265 87.310 ;
        RECT 31.455 87.140 31.625 87.310 ;
        RECT 34.125 87.140 34.295 87.310 ;
        RECT 34.485 87.140 34.655 87.310 ;
        RECT 36.855 87.140 37.025 87.310 ;
        RECT 37.215 87.140 37.385 87.310 ;
        RECT 39.885 87.140 40.055 87.310 ;
        RECT 40.245 87.140 40.415 87.310 ;
        RECT 42.615 87.140 42.785 87.310 ;
        RECT 42.975 87.140 43.145 87.310 ;
        RECT 45.645 87.140 45.815 87.310 ;
        RECT 46.005 87.140 46.175 87.310 ;
        RECT 48.375 87.140 48.545 87.310 ;
        RECT 48.735 87.140 48.905 87.310 ;
        RECT 52.930 87.185 53.100 87.355 ;
        RECT 53.410 87.185 53.580 87.355 ;
        RECT 53.880 87.185 54.050 87.355 ;
        RECT 54.360 87.185 54.530 87.355 ;
        RECT 54.900 87.185 55.070 87.355 ;
        RECT 55.380 87.185 55.550 87.355 ;
        RECT 55.855 87.185 56.025 87.355 ;
        RECT 56.335 87.185 56.505 87.355 ;
        RECT 56.895 87.185 57.065 87.355 ;
        RECT 57.375 87.185 57.545 87.355 ;
        RECT 57.850 87.185 58.020 87.355 ;
        RECT 58.330 87.185 58.500 87.355 ;
        RECT 58.870 87.185 59.040 87.355 ;
        RECT 59.350 87.185 59.520 87.355 ;
        RECT 59.825 87.185 59.995 87.355 ;
        RECT 60.305 87.185 60.475 87.355 ;
        RECT 60.895 87.185 61.065 87.355 ;
        RECT 61.375 87.185 61.545 87.355 ;
        RECT 61.850 87.185 62.020 87.355 ;
        RECT 62.330 87.185 62.500 87.355 ;
        RECT 62.870 87.185 63.040 87.355 ;
        RECT 63.350 87.185 63.520 87.355 ;
        RECT 63.825 87.185 63.995 87.355 ;
        RECT 64.305 87.185 64.475 87.355 ;
        RECT 64.865 87.185 65.035 87.355 ;
        RECT 65.345 87.185 65.515 87.355 ;
        RECT 65.820 87.185 65.990 87.355 ;
        RECT 66.300 87.185 66.470 87.355 ;
        RECT 66.840 87.185 67.010 87.355 ;
        RECT 67.320 87.185 67.490 87.355 ;
        RECT 67.795 87.185 67.965 87.355 ;
        RECT 68.275 87.185 68.445 87.355 ;
        RECT 52.930 86.825 53.100 86.995 ;
        RECT 53.410 86.825 53.580 86.995 ;
        RECT 53.880 86.825 54.050 86.995 ;
        RECT 54.360 86.825 54.530 86.995 ;
        RECT 54.900 86.825 55.070 86.995 ;
        RECT 55.380 86.825 55.550 86.995 ;
        RECT 55.855 86.825 56.025 86.995 ;
        RECT 56.335 86.825 56.505 86.995 ;
        RECT 56.895 86.825 57.065 86.995 ;
        RECT 57.375 86.825 57.545 86.995 ;
        RECT 57.850 86.825 58.020 86.995 ;
        RECT 58.330 86.825 58.500 86.995 ;
        RECT 58.870 86.825 59.040 86.995 ;
        RECT 59.350 86.825 59.520 86.995 ;
        RECT 59.825 86.825 59.995 86.995 ;
        RECT 60.305 86.825 60.475 86.995 ;
        RECT 60.895 86.825 61.065 86.995 ;
        RECT 61.375 86.825 61.545 86.995 ;
        RECT 61.850 86.825 62.020 86.995 ;
        RECT 62.330 86.825 62.500 86.995 ;
        RECT 62.870 86.825 63.040 86.995 ;
        RECT 63.350 86.825 63.520 86.995 ;
        RECT 63.825 86.825 63.995 86.995 ;
        RECT 64.305 86.825 64.475 86.995 ;
        RECT 64.865 86.825 65.035 86.995 ;
        RECT 65.345 86.825 65.515 86.995 ;
        RECT 65.820 86.825 65.990 86.995 ;
        RECT 66.300 86.825 66.470 86.995 ;
        RECT 66.840 86.825 67.010 86.995 ;
        RECT 67.320 86.825 67.490 86.995 ;
        RECT 67.795 86.825 67.965 86.995 ;
        RECT 68.275 86.825 68.445 86.995 ;
        RECT 16.845 86.060 17.015 86.230 ;
        RECT 17.205 86.060 17.375 86.230 ;
        RECT 19.575 86.060 19.745 86.230 ;
        RECT 19.935 86.060 20.105 86.230 ;
        RECT 22.605 86.060 22.775 86.230 ;
        RECT 22.965 86.060 23.135 86.230 ;
        RECT 25.335 86.060 25.505 86.230 ;
        RECT 25.695 86.060 25.865 86.230 ;
        RECT 28.365 86.060 28.535 86.230 ;
        RECT 28.725 86.060 28.895 86.230 ;
        RECT 31.095 86.060 31.265 86.230 ;
        RECT 31.455 86.060 31.625 86.230 ;
        RECT 34.125 86.060 34.295 86.230 ;
        RECT 34.485 86.060 34.655 86.230 ;
        RECT 36.855 86.060 37.025 86.230 ;
        RECT 37.215 86.060 37.385 86.230 ;
        RECT 39.885 86.060 40.055 86.230 ;
        RECT 40.245 86.060 40.415 86.230 ;
        RECT 42.615 86.060 42.785 86.230 ;
        RECT 42.975 86.060 43.145 86.230 ;
        RECT 45.645 86.060 45.815 86.230 ;
        RECT 46.005 86.060 46.175 86.230 ;
        RECT 48.375 86.060 48.545 86.230 ;
        RECT 48.735 86.060 48.905 86.230 ;
        RECT 16.190 40.225 16.360 40.395 ;
        RECT 17.025 40.225 17.195 40.395 ;
        RECT 17.885 40.225 18.055 40.395 ;
        RECT 18.720 40.225 18.890 40.395 ;
        RECT 19.970 40.220 20.140 40.390 ;
        RECT 20.330 40.220 20.500 40.390 ;
        RECT 20.690 40.220 20.860 40.390 ;
        RECT 26.380 40.200 26.550 40.370 ;
        RECT 26.740 40.200 26.910 40.370 ;
        RECT 27.100 40.200 27.270 40.370 ;
        RECT 23.735 39.500 23.905 39.670 ;
        RECT 24.105 39.500 24.275 39.670 ;
        RECT 24.700 39.500 24.870 39.670 ;
        RECT 30.525 40.230 30.695 40.400 ;
        RECT 30.895 40.230 31.065 40.400 ;
        RECT 31.255 40.230 31.425 40.400 ;
        RECT 32.470 40.220 32.640 40.390 ;
        RECT 33.305 40.220 33.475 40.390 ;
        RECT 34.140 40.220 34.310 40.390 ;
        RECT 35.000 40.220 35.170 40.390 ;
        RECT 38.740 40.220 38.910 40.390 ;
        RECT 39.100 40.220 39.270 40.390 ;
        RECT 39.460 40.220 39.630 40.390 ;
        RECT 41.025 40.215 41.195 40.385 ;
        RECT 41.860 40.215 42.030 40.385 ;
        RECT 42.695 40.215 42.865 40.385 ;
        RECT 43.555 40.215 43.725 40.385 ;
        RECT 45.240 40.200 45.410 40.370 ;
        RECT 45.600 40.200 45.770 40.370 ;
        RECT 45.960 40.200 46.130 40.370 ;
        RECT 49.385 40.230 49.555 40.400 ;
        RECT 49.755 40.230 49.925 40.400 ;
        RECT 50.115 40.230 50.285 40.400 ;
        RECT 51.330 40.220 51.500 40.390 ;
        RECT 52.165 40.220 52.335 40.390 ;
        RECT 53.000 40.220 53.170 40.390 ;
        RECT 53.860 40.220 54.030 40.390 ;
        RECT 57.600 40.220 57.770 40.390 ;
        RECT 57.960 40.220 58.130 40.390 ;
        RECT 58.320 40.220 58.490 40.390 ;
        RECT 59.620 40.215 59.790 40.385 ;
        RECT 60.455 40.215 60.625 40.385 ;
        RECT 61.290 40.215 61.460 40.385 ;
        RECT 62.150 40.215 62.320 40.385 ;
        RECT 73.660 33.160 73.830 33.330 ;
        RECT 74.130 33.160 74.300 33.330 ;
        RECT 73.660 32.800 73.830 32.970 ;
        RECT 74.130 32.800 74.300 32.970 ;
        RECT 30.365 29.875 30.535 30.045 ;
        RECT 30.725 29.875 30.895 30.045 ;
        RECT 31.095 29.875 31.265 30.045 ;
        RECT 14.235 29.155 14.405 29.325 ;
        RECT 14.595 29.155 14.765 29.325 ;
        RECT 14.965 29.155 15.135 29.325 ;
        RECT 18.105 29.155 18.275 29.325 ;
        RECT 18.465 29.155 18.635 29.325 ;
        RECT 20.170 29.155 20.340 29.325 ;
        RECT 20.530 29.155 20.700 29.325 ;
        RECT 20.900 29.155 21.070 29.325 ;
        RECT 24.595 29.175 24.765 29.345 ;
        RECT 24.955 29.175 25.125 29.345 ;
        RECT 34.485 29.845 34.655 30.015 ;
        RECT 34.845 29.845 35.015 30.015 ;
        RECT 35.215 29.845 35.385 30.015 ;
        RECT 44.535 29.875 44.705 30.045 ;
        RECT 44.985 29.875 45.155 30.045 ;
        RECT 45.355 29.875 45.525 30.045 ;
        RECT 48.745 29.845 48.915 30.015 ;
        RECT 49.105 29.845 49.275 30.015 ;
        RECT 49.475 29.845 49.645 30.015 ;
        RECT 36.525 29.155 36.695 29.325 ;
        RECT 36.885 29.155 37.055 29.325 ;
        RECT 37.255 29.155 37.425 29.325 ;
        RECT 50.845 29.155 51.015 29.325 ;
        RECT 51.205 29.155 51.375 29.325 ;
        RECT 51.565 29.155 51.735 29.325 ;
        RECT 56.960 29.065 57.130 29.235 ;
        RECT 57.320 29.065 57.490 29.235 ;
        RECT 58.520 29.065 58.690 29.235 ;
        RECT 58.880 29.065 59.050 29.235 ;
        RECT 60.080 29.065 60.250 29.235 ;
        RECT 60.440 29.065 60.610 29.235 ;
        RECT 61.640 29.065 61.810 29.235 ;
        RECT 62.000 29.065 62.170 29.235 ;
        RECT 63.200 29.065 63.370 29.235 ;
        RECT 63.560 29.065 63.730 29.235 ;
        RECT 64.760 29.065 64.930 29.235 ;
        RECT 65.120 29.065 65.290 29.235 ;
        RECT 66.320 29.065 66.490 29.235 ;
        RECT 66.680 29.065 66.850 29.235 ;
        RECT 67.750 29.065 67.920 29.235 ;
        RECT 68.110 29.065 68.280 29.235 ;
        RECT 71.870 29.090 72.040 29.260 ;
        RECT 72.230 29.090 72.400 29.260 ;
      LAYER met1 ;
        RECT 16.315 119.435 21.025 120.635 ;
        RECT 23.345 119.435 30.660 120.635 ;
        RECT 33.160 119.435 50.500 120.635 ;
        RECT 54.900 117.435 59.310 118.730 ;
        RECT 62.830 117.435 69.610 118.730 ;
        RECT 54.900 110.705 59.310 111.985 ;
        RECT 62.830 110.705 69.610 111.985 ;
        RECT 16.315 107.530 21.030 108.710 ;
        RECT 23.345 107.530 30.665 108.710 ;
        RECT 33.160 107.530 50.505 108.710 ;
        RECT 20.100 104.485 23.790 104.960 ;
        RECT 24.780 104.485 25.070 104.515 ;
        RECT 26.340 104.485 26.630 104.515 ;
        RECT 27.900 104.485 28.190 104.515 ;
        RECT 29.460 104.485 29.750 104.515 ;
        RECT 31.020 104.485 31.310 104.515 ;
        RECT 20.100 104.315 31.310 104.485 ;
        RECT 20.100 104.285 23.790 104.315 ;
        RECT 24.780 104.285 25.070 104.315 ;
        RECT 26.340 104.285 26.630 104.315 ;
        RECT 27.900 104.285 28.190 104.315 ;
        RECT 29.460 104.285 29.750 104.315 ;
        RECT 31.020 104.285 31.310 104.315 ;
        RECT 37.380 104.485 41.070 104.960 ;
        RECT 42.060 104.485 42.350 104.515 ;
        RECT 43.620 104.485 43.910 104.515 ;
        RECT 45.180 104.485 45.470 104.515 ;
        RECT 46.740 104.485 47.030 104.515 ;
        RECT 48.300 104.485 48.590 104.515 ;
        RECT 37.380 104.315 48.590 104.485 ;
        RECT 37.380 104.285 41.070 104.315 ;
        RECT 42.060 104.285 42.350 104.315 ;
        RECT 43.620 104.285 43.910 104.315 ;
        RECT 45.180 104.285 45.470 104.315 ;
        RECT 46.740 104.285 47.030 104.315 ;
        RECT 48.300 104.285 48.590 104.315 ;
        RECT 54.660 104.485 54.950 104.515 ;
        RECT 56.220 104.485 56.510 104.515 ;
        RECT 57.780 104.485 58.070 104.515 ;
        RECT 59.340 104.485 59.630 104.515 ;
        RECT 60.900 104.485 61.190 104.515 ;
        RECT 62.400 104.485 69.615 104.960 ;
        RECT 54.660 104.315 69.615 104.485 ;
        RECT 54.660 104.285 54.950 104.315 ;
        RECT 56.220 104.285 56.510 104.315 ;
        RECT 57.780 104.285 58.070 104.315 ;
        RECT 59.340 104.285 59.630 104.315 ;
        RECT 60.900 104.285 61.190 104.315 ;
        RECT 62.400 104.285 69.615 104.315 ;
        RECT 15.555 103.400 16.505 103.950 ;
        RECT 18.360 103.820 20.165 103.970 ;
        RECT 18.360 103.745 21.755 103.820 ;
        RECT 22.260 103.745 22.910 103.775 ;
        RECT 23.820 103.745 24.470 103.775 ;
        RECT 25.380 103.745 26.030 103.775 ;
        RECT 26.940 103.745 27.590 103.775 ;
        RECT 28.500 103.745 29.150 103.775 ;
        RECT 30.060 103.745 30.710 103.775 ;
        RECT 18.360 103.630 30.710 103.745 ;
        RECT 19.825 103.575 30.710 103.630 ;
        RECT 19.825 103.480 21.755 103.575 ;
        RECT 22.260 103.545 22.910 103.575 ;
        RECT 23.820 103.545 24.470 103.575 ;
        RECT 25.380 103.545 26.030 103.575 ;
        RECT 26.940 103.545 27.590 103.575 ;
        RECT 28.500 103.545 29.150 103.575 ;
        RECT 30.060 103.545 30.710 103.575 ;
        RECT 32.655 103.400 33.605 103.950 ;
        RECT 35.640 103.820 37.445 103.970 ;
        RECT 35.640 103.745 39.035 103.820 ;
        RECT 39.540 103.745 40.190 103.775 ;
        RECT 41.100 103.745 41.750 103.775 ;
        RECT 42.660 103.745 43.310 103.775 ;
        RECT 44.220 103.745 44.870 103.775 ;
        RECT 45.780 103.745 46.430 103.775 ;
        RECT 47.340 103.745 47.990 103.775 ;
        RECT 35.640 103.630 47.990 103.745 ;
        RECT 37.105 103.575 47.990 103.630 ;
        RECT 37.105 103.480 39.035 103.575 ;
        RECT 39.540 103.545 40.190 103.575 ;
        RECT 41.100 103.545 41.750 103.575 ;
        RECT 42.660 103.545 43.310 103.575 ;
        RECT 44.220 103.545 44.870 103.575 ;
        RECT 45.780 103.545 46.430 103.575 ;
        RECT 47.340 103.545 47.990 103.575 ;
        RECT 50.085 103.400 51.035 103.950 ;
        RECT 52.910 103.820 54.715 103.970 ;
        RECT 52.910 103.745 56.305 103.820 ;
        RECT 56.820 103.745 57.470 103.775 ;
        RECT 58.380 103.745 59.030 103.775 ;
        RECT 59.940 103.745 60.590 103.775 ;
        RECT 61.500 103.745 62.150 103.775 ;
        RECT 63.060 103.745 63.710 103.775 ;
        RECT 64.620 103.745 65.270 103.775 ;
        RECT 52.910 103.630 65.270 103.745 ;
        RECT 54.375 103.575 65.270 103.630 ;
        RECT 54.375 103.480 56.305 103.575 ;
        RECT 56.820 103.545 57.470 103.575 ;
        RECT 58.380 103.545 59.030 103.575 ;
        RECT 59.940 103.545 60.590 103.575 ;
        RECT 61.500 103.545 62.150 103.575 ;
        RECT 63.060 103.545 63.710 103.575 ;
        RECT 64.620 103.545 65.270 103.575 ;
        RECT 15.555 100.070 16.505 100.620 ;
        RECT 19.825 100.415 21.795 100.555 ;
        RECT 22.260 100.415 22.910 100.445 ;
        RECT 23.820 100.415 24.470 100.445 ;
        RECT 25.380 100.415 26.030 100.445 ;
        RECT 26.940 100.415 27.590 100.445 ;
        RECT 28.500 100.415 29.150 100.445 ;
        RECT 30.060 100.415 30.710 100.445 ;
        RECT 19.825 100.350 30.710 100.415 ;
        RECT 18.360 100.245 30.710 100.350 ;
        RECT 18.360 100.215 21.795 100.245 ;
        RECT 22.260 100.215 22.910 100.245 ;
        RECT 23.820 100.215 24.470 100.245 ;
        RECT 25.380 100.215 26.030 100.245 ;
        RECT 26.940 100.215 27.590 100.245 ;
        RECT 28.500 100.215 29.150 100.245 ;
        RECT 30.060 100.215 30.710 100.245 ;
        RECT 18.360 100.010 20.165 100.215 ;
        RECT 32.810 100.070 33.760 100.620 ;
        RECT 37.105 100.415 38.975 100.555 ;
        RECT 39.540 100.415 40.190 100.445 ;
        RECT 41.100 100.415 41.750 100.445 ;
        RECT 42.660 100.415 43.310 100.445 ;
        RECT 44.220 100.415 44.870 100.445 ;
        RECT 45.780 100.415 46.430 100.445 ;
        RECT 47.340 100.415 47.990 100.445 ;
        RECT 37.105 100.355 47.990 100.415 ;
        RECT 35.640 100.245 47.990 100.355 ;
        RECT 35.640 100.215 38.975 100.245 ;
        RECT 39.540 100.215 40.190 100.245 ;
        RECT 41.100 100.215 41.750 100.245 ;
        RECT 42.660 100.215 43.310 100.245 ;
        RECT 44.220 100.215 44.870 100.245 ;
        RECT 45.780 100.215 46.430 100.245 ;
        RECT 47.340 100.215 47.990 100.245 ;
        RECT 35.640 100.015 37.445 100.215 ;
        RECT 50.100 100.070 51.050 100.620 ;
        RECT 54.375 100.415 56.205 100.555 ;
        RECT 56.820 100.415 57.470 100.445 ;
        RECT 58.380 100.415 59.030 100.445 ;
        RECT 59.940 100.415 60.590 100.445 ;
        RECT 61.500 100.415 62.150 100.445 ;
        RECT 63.060 100.415 63.710 100.445 ;
        RECT 64.620 100.415 65.270 100.445 ;
        RECT 54.375 100.370 65.270 100.415 ;
        RECT 52.910 100.245 65.270 100.370 ;
        RECT 52.910 100.215 56.205 100.245 ;
        RECT 56.820 100.215 57.470 100.245 ;
        RECT 58.380 100.215 59.030 100.245 ;
        RECT 59.940 100.215 60.590 100.245 ;
        RECT 61.500 100.215 62.150 100.245 ;
        RECT 63.060 100.215 63.710 100.245 ;
        RECT 64.620 100.215 65.270 100.245 ;
        RECT 52.910 100.030 54.715 100.215 ;
        RECT 20.100 99.675 24.270 99.705 ;
        RECT 24.780 99.675 25.070 99.705 ;
        RECT 26.340 99.675 26.630 99.705 ;
        RECT 27.900 99.675 28.190 99.705 ;
        RECT 29.460 99.675 29.750 99.705 ;
        RECT 31.020 99.675 31.310 99.705 ;
        RECT 20.100 99.505 31.310 99.675 ;
        RECT 20.100 99.030 24.270 99.505 ;
        RECT 24.780 99.475 25.070 99.505 ;
        RECT 26.340 99.475 26.630 99.505 ;
        RECT 27.900 99.475 28.190 99.505 ;
        RECT 29.460 99.475 29.750 99.505 ;
        RECT 31.020 99.475 31.310 99.505 ;
        RECT 37.380 99.675 41.550 99.705 ;
        RECT 42.060 99.675 42.350 99.705 ;
        RECT 43.620 99.675 43.910 99.705 ;
        RECT 45.180 99.675 45.470 99.705 ;
        RECT 46.740 99.675 47.030 99.705 ;
        RECT 48.300 99.675 48.590 99.705 ;
        RECT 37.380 99.505 48.590 99.675 ;
        RECT 37.380 99.030 41.550 99.505 ;
        RECT 42.060 99.475 42.350 99.505 ;
        RECT 43.620 99.475 43.910 99.505 ;
        RECT 45.180 99.475 45.470 99.505 ;
        RECT 46.740 99.475 47.030 99.505 ;
        RECT 48.300 99.475 48.590 99.505 ;
        RECT 53.215 99.675 57.385 99.705 ;
        RECT 57.780 99.675 58.070 99.705 ;
        RECT 59.340 99.675 59.630 99.705 ;
        RECT 60.900 99.675 61.190 99.705 ;
        RECT 62.460 99.675 62.750 99.705 ;
        RECT 64.020 99.675 64.310 99.705 ;
        RECT 65.580 99.675 65.870 99.705 ;
        RECT 53.215 99.505 65.870 99.675 ;
        RECT 53.215 99.030 57.385 99.505 ;
        RECT 57.780 99.475 58.070 99.505 ;
        RECT 59.340 99.475 59.630 99.505 ;
        RECT 60.900 99.475 61.190 99.505 ;
        RECT 62.460 99.475 62.750 99.505 ;
        RECT 64.020 99.475 64.310 99.505 ;
        RECT 65.580 99.475 65.870 99.505 ;
        RECT 16.705 95.960 17.435 96.150 ;
        RECT 19.515 95.960 20.270 96.150 ;
        RECT 16.705 95.670 20.270 95.960 ;
        RECT 22.465 95.960 23.195 96.150 ;
        RECT 25.275 95.960 26.030 96.150 ;
        RECT 22.465 95.670 26.030 95.960 ;
        RECT 28.225 95.960 28.955 96.150 ;
        RECT 31.035 95.960 31.790 96.150 ;
        RECT 28.225 95.670 31.790 95.960 ;
        RECT 33.985 95.960 34.715 96.150 ;
        RECT 36.795 95.960 37.550 96.150 ;
        RECT 33.985 95.670 37.550 95.960 ;
        RECT 39.745 95.960 40.475 96.150 ;
        RECT 42.555 95.960 43.310 96.150 ;
        RECT 39.745 95.670 43.310 95.960 ;
        RECT 45.505 95.960 46.235 96.150 ;
        RECT 48.315 95.960 49.070 96.150 ;
        RECT 45.505 95.670 49.070 95.960 ;
        RECT 16.695 91.725 17.425 95.360 ;
        RECT 17.740 92.065 18.915 94.945 ;
        RECT 19.315 91.660 20.280 95.360 ;
        RECT 22.455 91.725 23.185 95.360 ;
        RECT 23.500 92.065 24.675 94.945 ;
        RECT 25.075 91.660 26.040 95.360 ;
        RECT 28.215 91.725 28.945 95.360 ;
        RECT 29.260 92.065 30.435 94.945 ;
        RECT 30.835 91.660 31.800 95.360 ;
        RECT 33.975 91.725 34.705 95.360 ;
        RECT 35.020 92.065 36.195 94.945 ;
        RECT 36.595 91.660 37.560 95.360 ;
        RECT 39.735 91.725 40.465 95.360 ;
        RECT 40.780 92.065 41.955 94.945 ;
        RECT 42.355 91.660 43.320 95.360 ;
        RECT 45.495 91.725 46.225 95.360 ;
        RECT 46.540 92.065 47.715 94.945 ;
        RECT 48.115 91.660 49.080 95.360 ;
        RECT 52.825 93.360 69.085 94.640 ;
        RECT 16.605 86.995 17.425 90.870 ;
        RECT 17.975 87.470 18.915 90.475 ;
        RECT 19.335 86.995 20.275 90.935 ;
        RECT 22.365 86.995 23.185 90.870 ;
        RECT 23.735 87.470 24.675 90.475 ;
        RECT 25.095 86.995 26.035 90.935 ;
        RECT 28.125 86.995 28.945 90.870 ;
        RECT 29.495 87.470 30.435 90.475 ;
        RECT 30.855 86.995 31.795 90.935 ;
        RECT 33.885 86.995 34.705 90.870 ;
        RECT 35.255 87.470 36.195 90.475 ;
        RECT 36.615 86.995 37.555 90.935 ;
        RECT 39.645 86.995 40.465 90.870 ;
        RECT 41.015 87.470 41.955 90.475 ;
        RECT 42.375 86.995 43.315 90.935 ;
        RECT 45.405 86.995 46.225 90.870 ;
        RECT 46.775 87.470 47.715 90.475 ;
        RECT 48.135 86.995 49.075 90.935 ;
        RECT 52.825 86.615 69.085 87.910 ;
        RECT 16.605 86.095 20.275 86.400 ;
        RECT 16.605 85.915 17.510 86.095 ;
        RECT 19.515 85.915 20.275 86.095 ;
        RECT 22.365 86.095 26.035 86.400 ;
        RECT 22.365 85.915 23.270 86.095 ;
        RECT 25.275 85.915 26.035 86.095 ;
        RECT 28.125 86.095 31.795 86.400 ;
        RECT 28.125 85.915 29.030 86.095 ;
        RECT 31.035 85.915 31.795 86.095 ;
        RECT 33.885 86.095 37.555 86.400 ;
        RECT 33.885 85.915 34.790 86.095 ;
        RECT 36.795 85.915 37.555 86.095 ;
        RECT 39.645 86.095 43.315 86.400 ;
        RECT 39.645 85.915 40.550 86.095 ;
        RECT 42.555 85.915 43.315 86.095 ;
        RECT 45.405 86.095 49.075 86.400 ;
        RECT 45.405 85.915 46.310 86.095 ;
        RECT 48.315 85.915 49.075 86.095 ;
        RECT 33.570 44.955 49.600 45.295 ;
        RECT 32.485 44.065 45.450 44.405 ;
        RECT 45.110 42.820 45.450 44.065 ;
        RECT 49.260 42.765 49.600 44.955 ;
        RECT 16.060 40.060 21.110 40.525 ;
        RECT 26.070 40.100 27.450 40.490 ;
        RECT 30.070 40.160 35.370 40.450 ;
        RECT 38.450 40.160 44.005 40.450 ;
        RECT 23.440 39.440 24.975 39.730 ;
        RECT 38.450 39.660 39.815 40.160 ;
        RECT 44.930 40.100 46.310 40.490 ;
        RECT 48.930 40.160 54.230 40.450 ;
        RECT 57.215 40.160 62.505 40.450 ;
        RECT 73.505 32.500 74.515 33.585 ;
        RECT 20.800 29.820 24.235 30.160 ;
        RECT 20.800 29.410 21.140 29.820 ;
        RECT 13.850 29.095 15.330 29.385 ;
        RECT 17.845 29.095 19.425 29.385 ;
        RECT 19.855 29.070 21.140 29.410 ;
        RECT 23.895 29.425 24.235 29.820 ;
        RECT 30.045 29.815 31.625 30.105 ;
        RECT 34.295 29.725 35.645 30.125 ;
        RECT 36.310 29.810 39.760 30.250 ;
        RECT 44.305 29.815 45.885 30.105 ;
        RECT 23.895 29.085 25.410 29.425 ;
        RECT 36.310 28.710 37.975 29.810 ;
        RECT 48.555 29.725 49.905 30.125 ;
        RECT 50.560 28.710 52.030 29.410 ;
        RECT 56.900 29.235 57.550 29.265 ;
        RECT 58.460 29.235 59.110 29.265 ;
        RECT 60.020 29.235 60.670 29.265 ;
        RECT 61.580 29.235 62.230 29.265 ;
        RECT 63.140 29.235 63.790 29.265 ;
        RECT 64.700 29.235 65.350 29.265 ;
        RECT 66.260 29.235 66.910 29.265 ;
        RECT 67.720 29.235 68.340 29.265 ;
        RECT 56.830 29.065 68.340 29.235 ;
        RECT 56.900 29.035 57.550 29.065 ;
        RECT 58.460 29.035 59.110 29.065 ;
        RECT 60.020 29.035 60.670 29.065 ;
        RECT 61.580 29.035 62.230 29.065 ;
        RECT 63.140 29.035 63.790 29.065 ;
        RECT 64.700 29.035 65.350 29.065 ;
        RECT 66.260 29.035 66.910 29.065 ;
        RECT 67.720 29.035 68.340 29.065 ;
        RECT 69.150 29.025 72.810 29.340 ;
        RECT 48.435 25.995 58.595 26.495 ;
      LAYER via ;
        RECT 17.655 119.795 17.915 120.055 ;
        RECT 17.995 119.795 18.255 120.055 ;
        RECT 18.315 119.795 18.575 120.055 ;
        RECT 18.720 119.795 18.980 120.055 ;
        RECT 19.060 119.795 19.320 120.055 ;
        RECT 19.380 119.795 19.640 120.055 ;
        RECT 24.355 119.865 24.615 120.125 ;
        RECT 24.695 119.865 24.955 120.125 ;
        RECT 25.015 119.865 25.275 120.125 ;
        RECT 25.420 119.865 25.680 120.125 ;
        RECT 25.760 119.865 26.020 120.125 ;
        RECT 26.080 119.865 26.340 120.125 ;
        RECT 34.275 119.940 34.535 120.200 ;
        RECT 34.615 119.940 34.875 120.200 ;
        RECT 34.935 119.940 35.195 120.200 ;
        RECT 35.340 119.940 35.600 120.200 ;
        RECT 35.680 119.940 35.940 120.200 ;
        RECT 36.000 119.940 36.260 120.200 ;
        RECT 36.485 119.940 36.745 120.200 ;
        RECT 36.825 119.940 37.085 120.200 ;
        RECT 55.485 117.915 55.745 118.175 ;
        RECT 55.825 117.915 56.085 118.175 ;
        RECT 56.145 117.915 56.405 118.175 ;
        RECT 67.645 117.900 67.905 118.160 ;
        RECT 67.985 117.900 68.245 118.160 ;
        RECT 68.305 117.900 68.565 118.160 ;
        RECT 55.085 111.170 55.345 111.430 ;
        RECT 55.425 111.170 55.685 111.430 ;
        RECT 55.745 111.170 56.005 111.430 ;
        RECT 56.150 111.170 56.410 111.430 ;
        RECT 56.490 111.170 56.750 111.430 ;
        RECT 56.810 111.170 57.070 111.430 ;
        RECT 68.410 111.005 68.670 111.265 ;
        RECT 68.750 111.005 69.010 111.265 ;
        RECT 69.070 111.005 69.330 111.265 ;
        RECT 17.185 108.060 17.445 108.320 ;
        RECT 17.525 108.060 17.785 108.320 ;
        RECT 17.845 108.060 18.105 108.320 ;
        RECT 18.250 108.060 18.510 108.320 ;
        RECT 18.590 108.060 18.850 108.320 ;
        RECT 18.910 108.060 19.170 108.320 ;
        RECT 23.915 107.940 24.175 108.200 ;
        RECT 24.255 107.940 24.515 108.200 ;
        RECT 24.575 107.940 24.835 108.200 ;
        RECT 24.980 107.940 25.240 108.200 ;
        RECT 25.320 107.940 25.580 108.200 ;
        RECT 25.640 107.940 25.900 108.200 ;
        RECT 34.275 107.955 34.535 108.215 ;
        RECT 34.615 107.955 34.875 108.215 ;
        RECT 34.935 107.955 35.195 108.215 ;
        RECT 35.340 107.955 35.600 108.215 ;
        RECT 35.680 107.955 35.940 108.215 ;
        RECT 36.000 107.955 36.260 108.215 ;
        RECT 36.485 107.955 36.745 108.215 ;
        RECT 36.825 107.955 37.085 108.215 ;
        RECT 20.305 104.615 20.565 104.875 ;
        RECT 20.645 104.615 20.905 104.875 ;
        RECT 20.965 104.615 21.225 104.875 ;
        RECT 21.370 104.615 21.630 104.875 ;
        RECT 21.710 104.615 21.970 104.875 ;
        RECT 22.030 104.615 22.290 104.875 ;
        RECT 22.515 104.615 22.775 104.875 ;
        RECT 22.855 104.615 23.115 104.875 ;
        RECT 37.585 104.615 37.845 104.875 ;
        RECT 37.925 104.615 38.185 104.875 ;
        RECT 38.245 104.615 38.505 104.875 ;
        RECT 38.650 104.615 38.910 104.875 ;
        RECT 38.990 104.615 39.250 104.875 ;
        RECT 39.310 104.615 39.570 104.875 ;
        RECT 39.795 104.615 40.055 104.875 ;
        RECT 40.135 104.615 40.395 104.875 ;
        RECT 66.925 104.570 67.185 104.830 ;
        RECT 67.265 104.570 67.525 104.830 ;
        RECT 67.585 104.570 67.845 104.830 ;
        RECT 67.990 104.570 68.250 104.830 ;
        RECT 68.330 104.570 68.590 104.830 ;
        RECT 15.660 103.530 15.920 103.790 ;
        RECT 16.000 103.530 16.260 103.790 ;
        RECT 32.760 103.530 33.020 103.790 ;
        RECT 33.100 103.530 33.360 103.790 ;
        RECT 50.190 103.530 50.450 103.790 ;
        RECT 50.530 103.530 50.790 103.790 ;
        RECT 15.660 100.200 15.920 100.460 ;
        RECT 16.000 100.200 16.260 100.460 ;
        RECT 32.915 100.200 33.175 100.460 ;
        RECT 33.255 100.200 33.515 100.460 ;
        RECT 50.205 100.200 50.465 100.460 ;
        RECT 50.545 100.200 50.805 100.460 ;
        RECT 21.045 99.110 21.305 99.370 ;
        RECT 21.385 99.110 21.645 99.370 ;
        RECT 21.705 99.110 21.965 99.370 ;
        RECT 22.215 99.110 22.475 99.370 ;
        RECT 22.555 99.110 22.815 99.370 ;
        RECT 22.875 99.110 23.135 99.370 ;
        RECT 37.860 99.075 38.120 99.335 ;
        RECT 38.200 99.075 38.460 99.335 ;
        RECT 38.520 99.075 38.780 99.335 ;
        RECT 39.030 99.075 39.290 99.335 ;
        RECT 39.370 99.075 39.630 99.335 ;
        RECT 39.690 99.075 39.950 99.335 ;
        RECT 53.695 99.400 53.955 99.660 ;
        RECT 54.035 99.400 54.295 99.660 ;
        RECT 54.355 99.400 54.615 99.660 ;
        RECT 54.865 99.400 55.125 99.660 ;
        RECT 55.205 99.400 55.465 99.660 ;
        RECT 55.525 99.400 55.785 99.660 ;
        RECT 18.540 95.690 18.800 95.950 ;
        RECT 18.860 95.690 19.120 95.950 ;
        RECT 24.300 95.690 24.560 95.950 ;
        RECT 24.620 95.690 24.880 95.950 ;
        RECT 30.060 95.690 30.320 95.950 ;
        RECT 30.380 95.690 30.640 95.950 ;
        RECT 35.820 95.690 36.080 95.950 ;
        RECT 36.140 95.690 36.400 95.950 ;
        RECT 41.580 95.690 41.840 95.950 ;
        RECT 41.900 95.690 42.160 95.950 ;
        RECT 47.340 95.690 47.600 95.950 ;
        RECT 47.660 95.690 47.920 95.950 ;
        RECT 17.805 94.460 18.065 94.720 ;
        RECT 17.805 94.140 18.065 94.400 ;
        RECT 17.805 93.800 18.065 94.060 ;
        RECT 17.805 93.480 18.065 93.740 ;
        RECT 17.805 93.140 18.065 93.400 ;
        RECT 17.805 92.800 18.065 93.060 ;
        RECT 19.730 93.950 19.990 94.210 ;
        RECT 19.730 93.625 19.990 93.885 ;
        RECT 19.730 93.295 19.990 93.555 ;
        RECT 19.730 92.900 19.990 93.160 ;
        RECT 19.730 92.575 19.990 92.835 ;
        RECT 19.730 92.245 19.990 92.505 ;
        RECT 22.720 94.885 22.980 95.145 ;
        RECT 22.720 94.560 22.980 94.820 ;
        RECT 22.720 94.230 22.980 94.490 ;
        RECT 22.720 93.835 22.980 94.095 ;
        RECT 22.720 93.510 22.980 93.770 ;
        RECT 22.720 93.180 22.980 93.440 ;
        RECT 23.565 94.460 23.825 94.720 ;
        RECT 23.565 94.140 23.825 94.400 ;
        RECT 23.565 93.800 23.825 94.060 ;
        RECT 23.565 93.480 23.825 93.740 ;
        RECT 23.565 93.140 23.825 93.400 ;
        RECT 23.565 92.800 23.825 93.060 ;
        RECT 28.435 94.255 28.695 94.515 ;
        RECT 28.435 93.930 28.695 94.190 ;
        RECT 28.435 93.600 28.695 93.860 ;
        RECT 28.435 93.205 28.695 93.465 ;
        RECT 28.435 92.880 28.695 93.140 ;
        RECT 28.435 92.550 28.695 92.810 ;
        RECT 29.325 94.460 29.585 94.720 ;
        RECT 29.325 94.140 29.585 94.400 ;
        RECT 29.325 93.800 29.585 94.060 ;
        RECT 29.325 93.480 29.585 93.740 ;
        RECT 29.325 93.140 29.585 93.400 ;
        RECT 29.325 92.800 29.585 93.060 ;
        RECT 34.310 93.045 34.570 93.305 ;
        RECT 34.310 92.650 34.570 92.910 ;
        RECT 34.310 92.325 34.570 92.585 ;
        RECT 34.310 91.995 34.570 92.255 ;
        RECT 35.085 94.460 35.345 94.720 ;
        RECT 35.085 94.140 35.345 94.400 ;
        RECT 35.085 93.800 35.345 94.060 ;
        RECT 35.085 93.480 35.345 93.740 ;
        RECT 35.085 93.140 35.345 93.400 ;
        RECT 35.085 92.800 35.345 93.060 ;
        RECT 39.965 94.255 40.225 94.515 ;
        RECT 39.965 93.930 40.225 94.190 ;
        RECT 39.965 93.600 40.225 93.860 ;
        RECT 39.965 93.205 40.225 93.465 ;
        RECT 39.965 92.880 40.225 93.140 ;
        RECT 39.965 92.550 40.225 92.810 ;
        RECT 40.845 94.460 41.105 94.720 ;
        RECT 40.845 94.140 41.105 94.400 ;
        RECT 40.845 93.800 41.105 94.060 ;
        RECT 40.845 93.480 41.105 93.740 ;
        RECT 40.845 93.140 41.105 93.400 ;
        RECT 40.845 92.800 41.105 93.060 ;
        RECT 45.740 94.255 46.000 94.515 ;
        RECT 45.740 93.930 46.000 94.190 ;
        RECT 45.740 93.600 46.000 93.860 ;
        RECT 45.740 93.205 46.000 93.465 ;
        RECT 45.740 92.880 46.000 93.140 ;
        RECT 45.740 92.550 46.000 92.810 ;
        RECT 46.605 94.460 46.865 94.720 ;
        RECT 46.605 94.140 46.865 94.400 ;
        RECT 46.605 93.800 46.865 94.060 ;
        RECT 46.605 93.480 46.865 93.740 ;
        RECT 46.605 93.140 46.865 93.400 ;
        RECT 46.605 92.800 46.865 93.060 ;
        RECT 53.150 94.000 53.410 94.260 ;
        RECT 53.490 94.000 53.750 94.260 ;
        RECT 53.810 94.000 54.070 94.260 ;
        RECT 54.215 94.000 54.475 94.260 ;
        RECT 53.150 93.615 53.410 93.875 ;
        RECT 53.490 93.615 53.750 93.875 ;
        RECT 53.810 93.615 54.070 93.875 ;
        RECT 54.215 93.615 54.475 93.875 ;
        RECT 16.915 89.990 17.175 90.250 ;
        RECT 16.915 89.665 17.175 89.925 ;
        RECT 16.915 89.335 17.175 89.595 ;
        RECT 16.915 88.940 17.175 89.200 ;
        RECT 16.915 88.615 17.175 88.875 ;
        RECT 16.915 88.285 17.175 88.545 ;
        RECT 18.550 89.720 18.810 89.980 ;
        RECT 18.550 89.400 18.810 89.660 ;
        RECT 18.550 89.060 18.810 89.320 ;
        RECT 18.550 88.740 18.810 89.000 ;
        RECT 18.550 88.400 18.810 88.660 ;
        RECT 18.550 88.080 18.810 88.340 ;
        RECT 24.310 89.720 24.570 89.980 ;
        RECT 24.310 89.400 24.570 89.660 ;
        RECT 24.310 89.060 24.570 89.320 ;
        RECT 24.310 88.740 24.570 89.000 ;
        RECT 24.310 88.400 24.570 88.660 ;
        RECT 24.310 88.080 24.570 88.340 ;
        RECT 25.430 89.345 25.690 89.605 ;
        RECT 25.430 89.020 25.690 89.280 ;
        RECT 25.430 88.690 25.690 88.950 ;
        RECT 25.430 88.295 25.690 88.555 ;
        RECT 25.430 87.970 25.690 88.230 ;
        RECT 25.430 87.640 25.690 87.900 ;
        RECT 30.070 89.720 30.330 89.980 ;
        RECT 30.070 89.400 30.330 89.660 ;
        RECT 30.070 89.060 30.330 89.320 ;
        RECT 30.070 88.740 30.330 89.000 ;
        RECT 30.070 88.400 30.330 88.660 ;
        RECT 30.070 88.080 30.330 88.340 ;
        RECT 31.210 89.345 31.470 89.605 ;
        RECT 31.210 89.020 31.470 89.280 ;
        RECT 31.210 88.690 31.470 88.950 ;
        RECT 31.210 88.295 31.470 88.555 ;
        RECT 31.210 87.970 31.470 88.230 ;
        RECT 31.210 87.640 31.470 87.900 ;
        RECT 35.830 89.720 36.090 89.980 ;
        RECT 35.830 89.400 36.090 89.660 ;
        RECT 35.830 89.060 36.090 89.320 ;
        RECT 35.830 88.740 36.090 89.000 ;
        RECT 35.830 88.400 36.090 88.660 ;
        RECT 35.830 88.080 36.090 88.340 ;
        RECT 36.930 89.345 37.190 89.605 ;
        RECT 36.930 89.020 37.190 89.280 ;
        RECT 36.930 88.690 37.190 88.950 ;
        RECT 36.930 88.295 37.190 88.555 ;
        RECT 36.930 87.970 37.190 88.230 ;
        RECT 36.930 87.640 37.190 87.900 ;
        RECT 41.590 89.720 41.850 89.980 ;
        RECT 41.590 89.400 41.850 89.660 ;
        RECT 41.590 89.060 41.850 89.320 ;
        RECT 41.590 88.740 41.850 89.000 ;
        RECT 41.590 88.400 41.850 88.660 ;
        RECT 41.590 88.080 41.850 88.340 ;
        RECT 42.680 89.345 42.940 89.605 ;
        RECT 42.680 89.020 42.940 89.280 ;
        RECT 42.680 88.690 42.940 88.950 ;
        RECT 42.680 88.295 42.940 88.555 ;
        RECT 42.680 87.970 42.940 88.230 ;
        RECT 42.680 87.640 42.940 87.900 ;
        RECT 47.350 89.720 47.610 89.980 ;
        RECT 47.350 89.400 47.610 89.660 ;
        RECT 47.350 89.060 47.610 89.320 ;
        RECT 47.350 88.740 47.610 89.000 ;
        RECT 47.350 88.400 47.610 88.660 ;
        RECT 47.350 88.080 47.610 88.340 ;
        RECT 48.435 89.345 48.695 89.605 ;
        RECT 48.435 89.020 48.695 89.280 ;
        RECT 48.435 88.690 48.695 88.950 ;
        RECT 48.435 88.295 48.695 88.555 ;
        RECT 48.435 87.970 48.695 88.230 ;
        RECT 48.435 87.640 48.695 87.900 ;
        RECT 53.650 87.125 53.910 87.385 ;
        RECT 53.990 87.125 54.250 87.385 ;
        RECT 54.310 87.125 54.570 87.385 ;
        RECT 54.715 87.125 54.975 87.385 ;
        RECT 55.055 87.125 55.315 87.385 ;
        RECT 55.375 87.125 55.635 87.385 ;
        RECT 17.920 86.115 18.180 86.375 ;
        RECT 18.240 86.115 18.500 86.375 ;
        RECT 23.680 86.115 23.940 86.375 ;
        RECT 24.000 86.115 24.260 86.375 ;
        RECT 29.440 86.115 29.700 86.375 ;
        RECT 29.760 86.115 30.020 86.375 ;
        RECT 35.200 86.115 35.460 86.375 ;
        RECT 35.520 86.115 35.780 86.375 ;
        RECT 40.960 86.115 41.220 86.375 ;
        RECT 41.280 86.115 41.540 86.375 ;
        RECT 46.720 86.115 46.980 86.375 ;
        RECT 47.040 86.115 47.300 86.375 ;
        RECT 33.650 44.995 33.910 45.255 ;
        RECT 33.970 44.995 34.230 45.255 ;
        RECT 34.375 44.995 34.635 45.255 ;
        RECT 34.695 44.995 34.955 45.255 ;
        RECT 32.710 44.105 32.970 44.365 ;
        RECT 33.030 44.105 33.290 44.365 ;
        RECT 33.435 44.105 33.695 44.365 ;
        RECT 33.755 44.105 34.015 44.365 ;
        RECT 45.155 43.250 45.415 43.510 ;
        RECT 45.155 42.910 45.415 43.170 ;
        RECT 49.305 43.215 49.565 43.475 ;
        RECT 49.305 42.875 49.565 43.135 ;
        RECT 17.535 40.165 17.795 40.425 ;
        RECT 17.875 40.165 18.135 40.425 ;
        RECT 26.130 40.175 26.390 40.435 ;
        RECT 26.470 40.175 26.730 40.435 ;
        RECT 30.265 40.175 30.525 40.435 ;
        RECT 30.605 40.175 30.865 40.435 ;
        RECT 44.990 40.175 45.250 40.435 ;
        RECT 45.330 40.175 45.590 40.435 ;
        RECT 49.125 40.175 49.385 40.435 ;
        RECT 49.465 40.175 49.725 40.435 ;
        RECT 57.575 40.175 57.835 40.435 ;
        RECT 57.895 40.175 58.155 40.435 ;
        RECT 58.235 40.175 58.495 40.435 ;
        RECT 24.300 39.450 24.560 39.710 ;
        RECT 24.640 39.450 24.900 39.710 ;
        RECT 39.015 39.695 39.275 39.955 ;
        RECT 39.335 39.695 39.595 39.955 ;
        RECT 73.735 33.265 73.995 33.525 ;
        RECT 74.065 33.265 74.325 33.525 ;
        RECT 73.735 32.925 73.995 33.185 ;
        RECT 74.065 32.925 74.325 33.185 ;
        RECT 73.735 32.605 73.995 32.865 ;
        RECT 74.065 32.605 74.325 32.865 ;
        RECT 14.535 29.105 14.795 29.365 ;
        RECT 14.875 29.105 15.135 29.365 ;
        RECT 18.630 29.105 18.890 29.365 ;
        RECT 18.970 29.105 19.230 29.365 ;
        RECT 30.830 29.830 31.090 30.090 ;
        RECT 31.170 29.830 31.430 30.090 ;
        RECT 34.965 29.830 35.225 30.090 ;
        RECT 35.305 29.830 35.565 30.090 ;
        RECT 39.015 29.915 39.275 30.175 ;
        RECT 39.355 29.915 39.615 30.175 ;
        RECT 45.090 29.830 45.350 30.090 ;
        RECT 45.430 29.830 45.690 30.090 ;
        RECT 49.225 29.830 49.485 30.090 ;
        RECT 49.565 29.830 49.825 30.090 ;
        RECT 50.705 28.790 50.965 29.050 ;
        RECT 51.045 28.790 51.305 29.050 ;
        RECT 51.365 28.790 51.625 29.050 ;
        RECT 51.705 28.790 51.965 29.050 ;
        RECT 71.835 29.045 72.095 29.305 ;
        RECT 72.175 29.045 72.435 29.305 ;
        RECT 50.705 26.115 50.965 26.375 ;
        RECT 51.045 26.115 51.305 26.375 ;
        RECT 51.365 26.115 51.625 26.375 ;
        RECT 51.705 26.115 51.965 26.375 ;
        RECT 57.170 26.105 57.430 26.365 ;
        RECT 57.510 26.105 57.770 26.365 ;
        RECT 57.830 26.105 58.090 26.365 ;
        RECT 58.170 26.105 58.430 26.365 ;
      LAYER met2 ;
        RECT 16.660 119.750 20.680 120.090 ;
        RECT 23.615 119.835 27.310 120.175 ;
        RECT 33.690 119.905 38.320 120.245 ;
        RECT 16.660 108.365 17.000 119.750 ;
        RECT 16.660 108.025 20.390 108.365 ;
        RECT 20.050 104.925 20.390 108.025 ;
        RECT 23.615 108.255 23.955 119.835 ;
        RECT 33.690 108.265 34.030 119.905 ;
        RECT 55.170 117.805 56.855 118.305 ;
        RECT 67.425 117.805 69.445 118.305 ;
        RECT 55.170 111.550 55.670 117.805 ;
        RECT 45.385 111.050 57.245 111.550 ;
        RECT 68.945 111.380 69.445 117.805 ;
        RECT 23.615 107.915 26.270 108.255 ;
        RECT 20.050 104.585 23.745 104.925 ;
        RECT 13.170 103.495 17.430 103.835 ;
        RECT 13.170 96.650 13.510 103.495 ;
        RECT 14.515 100.185 17.795 100.525 ;
        RECT 14.515 97.840 14.855 100.185 ;
        RECT 25.930 99.420 26.270 107.915 ;
        RECT 33.470 107.925 39.350 108.265 ;
        RECT 33.470 104.925 33.810 107.925 ;
        RECT 33.470 104.585 41.235 104.925 ;
        RECT 20.755 99.080 26.270 99.420 ;
        RECT 29.275 103.485 34.935 103.825 ;
        RECT 14.515 97.500 23.885 97.840 ;
        RECT 13.170 96.310 18.120 96.650 ;
        RECT 17.780 94.775 18.120 96.310 ;
        RECT 18.445 95.635 19.210 95.995 ;
        RECT 16.890 43.595 17.230 90.490 ;
        RECT 17.740 86.375 18.145 94.775 ;
        RECT 18.445 87.980 18.885 95.635 ;
        RECT 17.740 86.095 18.575 86.375 ;
        RECT 19.695 44.535 20.035 94.595 ;
        RECT 22.675 48.505 23.015 95.215 ;
        RECT 23.545 94.775 23.885 97.500 ;
        RECT 24.205 95.635 24.970 95.995 ;
        RECT 23.500 86.375 23.905 94.775 ;
        RECT 24.205 87.980 24.645 95.635 ;
        RECT 29.275 94.775 29.615 103.485 ;
        RECT 32.600 100.165 35.365 100.505 ;
        RECT 29.965 95.635 30.730 95.995 ;
        RECT 23.500 86.095 24.335 86.375 ;
        RECT 25.390 49.755 25.730 89.750 ;
        RECT 28.380 51.245 28.720 94.750 ;
        RECT 29.260 86.375 29.665 94.775 ;
        RECT 29.965 87.980 30.405 95.635 ;
        RECT 35.025 94.775 35.365 100.165 ;
        RECT 45.385 99.450 45.885 111.050 ;
        RECT 68.290 110.880 69.445 111.380 ;
        RECT 68.290 104.960 68.790 110.880 ;
        RECT 66.780 104.460 68.790 104.960 ;
        RECT 37.275 98.950 45.885 99.450 ;
        RECT 47.835 103.490 51.035 103.830 ;
        RECT 47.835 98.160 48.175 103.490 ;
        RECT 49.975 100.135 52.530 100.475 ;
        RECT 40.800 97.820 48.175 98.160 ;
        RECT 35.725 95.635 36.490 95.995 ;
        RECT 29.260 86.095 30.095 86.375 ;
        RECT 31.160 53.090 31.500 90.440 ;
        RECT 34.260 54.850 34.600 93.415 ;
        RECT 35.020 86.375 35.425 94.775 ;
        RECT 35.725 87.980 36.165 95.635 ;
        RECT 35.020 86.095 35.855 86.375 ;
        RECT 36.885 56.290 37.225 90.590 ;
        RECT 36.885 55.950 37.670 56.290 ;
        RECT 34.260 54.510 36.430 54.850 ;
        RECT 31.160 52.750 33.895 53.090 ;
        RECT 28.380 50.905 32.195 51.245 ;
        RECT 25.390 49.415 30.730 49.755 ;
        RECT 22.675 48.165 26.570 48.505 ;
        RECT 19.695 44.195 24.770 44.535 ;
        RECT 16.890 43.255 18.015 43.595 ;
        RECT 17.675 40.520 18.015 43.255 ;
        RECT 17.400 40.060 18.220 40.520 ;
        RECT 24.430 39.930 24.770 44.195 ;
        RECT 26.230 40.635 26.570 48.165 ;
        RECT 26.025 40.060 26.870 40.635 ;
        RECT 30.390 40.600 30.730 49.415 ;
        RECT 31.855 44.405 32.195 50.905 ;
        RECT 33.555 45.295 33.895 52.750 ;
        RECT 33.555 44.955 35.065 45.295 ;
        RECT 31.855 44.065 34.190 44.405 ;
        RECT 36.090 43.090 36.430 54.510 ;
        RECT 34.775 42.750 36.430 43.090 ;
        RECT 30.160 40.060 31.000 40.600 ;
        RECT 24.180 39.300 24.975 39.930 ;
        RECT 34.775 33.630 35.115 42.750 ;
        RECT 37.330 42.020 37.670 55.950 ;
        RECT 14.505 33.290 35.115 33.630 ;
        RECT 35.960 41.680 37.670 42.020 ;
        RECT 14.505 29.460 14.845 33.290 ;
        RECT 35.960 32.890 36.300 41.680 ;
        RECT 39.920 41.195 40.260 94.970 ;
        RECT 40.800 94.775 41.140 97.820 ;
        RECT 52.190 97.130 52.530 100.135 ;
        RECT 46.560 96.790 52.530 97.130 ;
        RECT 53.525 99.360 55.945 99.700 ;
        RECT 41.485 95.635 42.250 95.995 ;
        RECT 40.780 86.375 41.185 94.775 ;
        RECT 41.485 87.980 41.925 95.635 ;
        RECT 46.560 94.775 46.900 96.790 ;
        RECT 47.245 95.635 48.010 95.995 ;
        RECT 40.780 86.095 41.615 86.375 ;
        RECT 18.750 32.550 36.300 32.890 ;
        RECT 36.765 40.855 40.260 41.195 ;
        RECT 14.440 28.955 15.210 29.460 ;
        RECT 18.750 29.450 19.090 32.550 ;
        RECT 36.765 32.115 37.105 40.855 ;
        RECT 42.645 40.645 42.985 90.655 ;
        RECT 45.690 48.650 46.030 94.600 ;
        RECT 46.540 86.375 46.945 94.775 ;
        RECT 47.245 87.980 47.685 95.635 ;
        RECT 53.525 94.330 53.865 99.360 ;
        RECT 52.980 93.535 54.770 94.330 ;
        RECT 46.540 86.095 47.375 86.375 ;
        RECT 48.390 50.645 48.730 90.915 ;
        RECT 53.525 87.425 53.865 93.535 ;
        RECT 53.525 87.085 55.940 87.425 ;
        RECT 48.390 50.305 55.795 50.645 ;
        RECT 45.690 48.310 53.180 48.650 ;
        RECT 30.985 31.775 37.105 32.115 ;
        RECT 37.545 40.305 42.985 40.645 ;
        RECT 45.110 40.590 45.450 43.565 ;
        RECT 30.985 30.225 31.325 31.775 ;
        RECT 37.545 31.095 37.885 40.305 ;
        RECT 44.885 40.060 45.730 40.590 ;
        RECT 49.260 40.540 49.600 43.615 ;
        RECT 49.020 40.060 49.860 40.540 ;
        RECT 35.095 30.755 37.885 31.095 ;
        RECT 35.095 30.235 35.435 30.755 ;
        RECT 30.705 29.715 31.535 30.225 ;
        RECT 34.840 29.715 35.670 30.235 ;
        RECT 38.935 29.890 39.740 39.970 ;
        RECT 52.840 33.420 53.180 48.310 ;
        RECT 45.170 33.080 53.180 33.420 ;
        RECT 45.170 30.220 45.510 33.080 ;
        RECT 55.455 32.405 55.795 50.305 ;
        RECT 49.380 32.065 55.795 32.405 ;
        RECT 49.380 30.260 49.720 32.065 ;
        RECT 44.965 29.715 45.795 30.220 ;
        RECT 49.100 29.715 49.930 30.260 ;
        RECT 18.495 28.955 19.305 29.450 ;
        RECT 14.505 28.935 14.845 28.955 ;
        RECT 50.625 25.905 52.035 29.165 ;
        RECT 57.165 25.940 58.565 40.560 ;
        RECT 73.415 32.380 74.640 33.745 ;
        RECT 73.875 29.350 74.215 32.380 ;
        RECT 71.750 29.010 74.215 29.350 ;
  END
END armleo_gpio
END LIBRARY

